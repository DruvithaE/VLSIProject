magic
tech scmos
timestamp 1698561877
<< nwell >>
rect -64 0 67 41
<< ntransistor >>
rect -38 -70 -31 -55
rect 26 -70 33 -55
<< ptransistor >>
rect -38 15 -31 30
rect 26 15 33 30
<< ndiffusion >>
rect -52 -57 -38 -55
rect -52 -64 -50 -57
rect -42 -64 -38 -57
rect -52 -70 -38 -64
rect -31 -58 -12 -55
rect -31 -67 -28 -58
rect -18 -67 -12 -58
rect -31 -70 -12 -67
rect 7 -56 26 -55
rect 7 -64 13 -56
rect 21 -64 26 -56
rect 7 -70 26 -64
rect 33 -57 47 -55
rect 33 -65 36 -57
rect 44 -65 47 -57
rect 33 -70 47 -65
<< pdiffusion >>
rect -52 28 -38 30
rect -52 22 -49 28
rect -42 22 -38 28
rect -52 15 -38 22
rect -31 26 -12 30
rect -31 18 -27 26
rect -18 18 -12 26
rect -31 15 -12 18
rect 15 26 26 30
rect 15 19 17 26
rect 25 19 26 26
rect 15 15 26 19
rect 33 24 55 30
rect 33 18 36 24
rect 44 18 55 24
rect 33 15 55 18
<< ndcontact >>
rect -50 -64 -42 -57
rect -28 -67 -18 -58
rect 13 -64 21 -56
rect 36 -65 44 -57
<< pdcontact >>
rect -49 22 -42 28
rect -27 18 -18 26
rect 17 19 25 26
rect 36 18 44 24
<< polysilicon >>
rect -38 30 -31 33
rect 26 30 33 33
rect -38 -55 -31 15
rect 26 -55 33 15
rect -38 -74 -31 -70
rect 26 -75 33 -70
<< metal1 >>
rect -49 42 25 48
rect -49 28 -42 42
rect 17 26 25 42
rect -27 -13 -18 18
rect 36 -13 44 18
rect -27 -21 44 -13
rect -28 -49 21 -41
rect -50 -86 -42 -64
rect -28 -58 -18 -49
rect 13 -56 21 -49
rect 36 -57 44 -21
<< labels >>
rlabel polysilicon -35 -19 -34 -15 1 x
rlabel polysilicon 28 -29 29 -25 1 y
rlabel metal1 -44 -82 -43 -78 1 gnd
rlabel metal1 -11 43 -10 47 5 vdd
rlabel metal1 39 -17 40 -13 1 out
<< end >>
