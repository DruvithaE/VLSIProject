
`include "mux.v"

module testbench;

    reg S0, S1;
    reg enable;
    reg [3:0] a, b;
    wire [4:0] Y;
    wire [3:0] y;
    wire Y4;

    assign y[3:0] = Y[3:0];
    assign Y4 = Y[4];

    mux inst1(.Y(Y),.S0(S0),.S1(S1),.a(a),.b(b),.enable(enable));
    initial begin
         #5   enable = 1;S0 =0;S1 =0; a = 4'b010;b = 4'b0001;
        $dumpfile("output.vcd"); 
        $dumpvars(S1,S1, S0, a[3:0], b[3:0], Y[4:0]);
        $monitor(" S1 =%b;S0 =%b; a = %b;b = %b; Y=%b; Y4=%b", S1 ,S0 ,a ,b ,Y[3:0],Y[4]);
        #5   a = 4'b0000; b = 4'b0000;
        #5   a = 4'b0000; b = 4'b0011;
        #5   a = 4'b0000; b = 4'b1111;
        #5 a = 4'b0001; b = 4'b0000;
        #5 a = 4'b0001; b = 4'b1100;
        #5 a = 4'b0001; b = 4'b1101;
        #5 a = 4'b0001; b = 4'b1111;
        #5 a = 4'b0010; b = 4'b0000;
        #5 a = 4'b0010; b = 4'b0001;
        #5 a = 4'b0010; b = 4'b0010;
        #5 a = 4'b0010; b = 4'b0100;
        #5 a = 4'b0010; b = 4'b0101;
        #5 a = 4'b0010; b = 4'b1110;
        #5 a = 4'b0010; b = 4'b1111;
        #5 a = 4'b0011; b = 4'b0000;
        #5 a = 4'b0011; b = 4'b0001;
        #5 a = 4'b0011; b = 4'b0010;
        #5 a = 4'b0011; b = 4'b0011;
        #5 a = 4'b0011; b = 4'b0100;
        #5 a = 4'b0011; b = 4'b0110;
        #5 a = 4'b0011; b = 4'b0111;
        #5 a = 4'b0011; b = 4'b1110;
        #5 a = 4'b0011; b = 4'b1111;
        #5 a = 4'b0100; b = 4'b0000;
        #5 a = 4'b0100; b = 4'b0001;
        #5 a = 4'b0100; b = 4'b0101;
        #5 a = 4'b0100; b = 4'b0111;
        #5 a = 4'b0100; b = 4'b1001;
        #5 a = 4'b0100; b = 4'b1010;
        #5 a = 4'b0100; b = 4'b1100;
        #5 a = 4'b0100; b = 4'b1110;
        #5 a = 4'b0101; b = 4'b0101;
        #5 a = 4'b0101; b = 4'b0110;
        #5 a = 4'b0101; b = 4'b0111;
        #5 a = 4'b0101; b = 4'b1001;
        #5 a = 4'b0101; b = 4'b1010;
        #5 a = 4'b0101; b = 4'b1101;
        #5 a = 4'b0101; b = 4'b1110;
        #5 a = 4'b0101; b = 4'b1111;
        #5 a = 4'b0110; b = 4'b0000;
        #5 a = 4'b0110; b = 4'b1101;
        #5 a = 4'b0110; b = 4'b1110;
        #5 a = 4'b0110; b = 4'b1111;
        #5 a = 4'b0111; b = 4'b0000;
        #5 a = 4'b0111; b = 4'b0010;
        #5 a = 4'b0111; b = 4'b0011;
        #5 a = 4'b0111; b = 4'b0111;
        #5 a = 4'b0111; b = 4'b1000;
        #5 a = 4'b0111; b = 4'b1101;
        #5 a = 4'b0111; b = 4'b1110;
        #5 a = 4'b1000; b = 4'b0000;
        #5 a = 4'b1000; b = 4'b0001;
        #5 a = 4'b1000; b = 4'b0010;
        #5 a = 4'b1000; b = 4'b1010;
        #5 a = 4'b1000; b = 4'b1100;
        #5 a = 4'b1000; b = 4'b1101;
        #5 a = 4'b1000; b = 4'b1111;
        #5 a = 4'b1110; b = 4'b0000;
        #5 a = 4'b1110; b = 4'b0011;
        #5 a = 4'b1110; b = 4'b0100;
        #5 a = 4'b1110; b = 4'b1001;
        #5 a = 4'b1110; b = 4'b1010;
        #5 a = 4'b1110; b = 4'b1011;
        #5 a = 4'b1110; b = 4'b1110;
        #5 a = 4'b1110; b = 4'b1111;
        #5 a = 4'b1101; b = 4'b0000;
        #5 a = 4'b1101; b = 4'b0001;
        #5 a = 4'b1101; b = 4'b0010;
        #5 a = 4'b1101; b = 4'b0110;
        #5 a = 4'b1101; b = 4'b0111;
        #5 a = 4'b1101; b = 4'b1010;
        #5 a = 4'b1101; b = 4'b1011;
        #5 a = 4'b1101; b = 4'b1100;
        #5 a = 4'b1101; b = 4'b1111;
        #5 a = 4'b1111; b = 4'b0000;
        #5 a = 4'b1111; b = 4'b0001;
        #5 a = 4'b1111; b = 4'b0010;
        #5 a = 4'b1111; b = 4'b0110;
        #5 a = 4'b1111; b = 4'b0111;
        #5 a = 4'b1111; b = 4'b1000;
        #5 a = 4'b1111; b = 4'b1001;
        #5 a = 4'b1111; b = 4'b1111;

        #5 $finish;
    end


endmodule

