magic
tech scmos
timestamp 1700152510
<< nwell >>
rect -989 724 -858 765
rect -786 724 -655 765
rect -599 724 -468 765
rect -418 724 -287 765
rect 105 445 236 486
rect 308 445 439 486
rect 495 445 626 486
rect 676 445 807 486
rect 845 439 976 480
rect 1048 439 1179 480
rect 1235 439 1366 480
rect 1416 439 1547 480
rect -961 377 -830 418
rect -758 377 -627 418
rect -571 377 -440 418
rect -390 377 -259 418
rect 5 153 136 194
rect 174 142 240 184
rect 288 149 419 190
rect 457 138 523 180
rect 552 153 640 178
rect 646 153 699 178
rect -961 -9 -830 32
rect -758 -9 -627 32
rect -571 -9 -440 32
rect -390 -9 -259 32
rect 162 -279 293 -238
rect 365 -279 496 -238
rect 552 -279 683 -238
rect 733 -279 864 -238
rect 902 -285 1033 -244
rect 1105 -285 1236 -244
rect 1292 -285 1423 -244
rect 1473 -285 1604 -244
rect -961 -433 -830 -392
rect -758 -433 -627 -392
rect -571 -433 -440 -392
rect -390 -433 -259 -392
rect 62 -571 193 -530
rect 231 -582 297 -540
rect 345 -575 476 -534
rect 514 -586 580 -544
rect 609 -571 697 -546
rect 703 -571 756 -546
rect 142 -869 273 -828
rect 345 -869 476 -828
rect 532 -869 663 -828
rect 713 -869 844 -828
rect 882 -875 1013 -834
rect 1085 -875 1216 -834
rect 1272 -875 1403 -834
rect 1453 -875 1584 -834
rect 42 -1161 173 -1120
rect 211 -1172 277 -1130
rect 325 -1165 456 -1124
rect 494 -1176 560 -1134
rect 589 -1161 677 -1136
rect 683 -1161 736 -1136
rect 170 -1493 301 -1452
rect 373 -1493 504 -1452
rect 560 -1493 691 -1452
rect 741 -1493 872 -1452
rect 910 -1499 1041 -1458
rect 1113 -1499 1244 -1458
rect 1300 -1499 1431 -1458
rect 1481 -1499 1612 -1458
rect 70 -1785 201 -1744
rect 239 -1796 305 -1754
rect 353 -1789 484 -1748
rect 522 -1800 588 -1758
rect 617 -1785 705 -1760
rect 711 -1785 764 -1760
<< ntransistor >>
rect -963 654 -956 669
rect -899 654 -892 669
rect -760 654 -753 669
rect -696 654 -689 669
rect -573 654 -566 669
rect -509 654 -502 669
rect -392 654 -385 669
rect -328 654 -321 669
rect -935 307 -928 322
rect -871 307 -864 322
rect -732 307 -725 322
rect -668 307 -661 322
rect -545 307 -538 322
rect -481 307 -474 322
rect -364 307 -357 322
rect -300 307 -293 322
rect -935 -79 -928 -64
rect -871 -79 -864 -64
rect -732 -79 -725 -64
rect -668 -79 -661 -64
rect -545 -79 -538 -64
rect -481 -79 -474 -64
rect -364 -79 -357 -64
rect -300 -79 -293 -64
rect -935 -503 -928 -488
rect -871 -503 -864 -488
rect -732 -503 -725 -488
rect -668 -503 -661 -488
rect -545 -503 -538 -488
rect -481 -503 -474 -488
rect -364 -503 -357 -488
rect -300 -503 -293 -488
rect 131 375 138 390
rect 195 375 202 390
rect 334 375 341 390
rect 398 375 405 390
rect 521 375 530 390
rect 585 375 592 390
rect 702 375 709 390
rect 766 375 773 390
rect 871 369 878 384
rect 935 369 942 384
rect 1074 369 1081 384
rect 1138 369 1145 384
rect 1261 369 1268 384
rect 1325 369 1332 384
rect 1442 369 1449 384
rect 1506 369 1513 384
rect 31 83 38 98
rect 95 83 102 98
rect 204 77 212 93
rect 314 79 321 94
rect 378 79 385 94
rect 574 99 580 110
rect 615 99 621 110
rect 666 99 672 110
rect 487 73 495 89
rect 188 -349 195 -334
rect 252 -349 259 -334
rect 391 -349 398 -334
rect 455 -349 462 -334
rect 578 -349 587 -334
rect 642 -349 649 -334
rect 759 -349 766 -334
rect 823 -349 830 -334
rect 928 -355 935 -340
rect 992 -355 999 -340
rect 1131 -355 1138 -340
rect 1195 -355 1202 -340
rect 1318 -355 1325 -340
rect 1382 -355 1389 -340
rect 1499 -355 1506 -340
rect 1563 -355 1570 -340
rect 88 -641 95 -626
rect 152 -641 159 -626
rect 261 -647 269 -631
rect 371 -645 378 -630
rect 435 -645 442 -630
rect 631 -625 637 -614
rect 672 -625 678 -614
rect 723 -625 729 -614
rect 544 -651 552 -635
rect 168 -939 175 -924
rect 232 -939 239 -924
rect 371 -939 378 -924
rect 435 -939 442 -924
rect 558 -939 567 -924
rect 622 -939 629 -924
rect 739 -939 746 -924
rect 803 -939 810 -924
rect 908 -945 915 -930
rect 972 -945 979 -930
rect 1111 -945 1118 -930
rect 1175 -945 1182 -930
rect 1298 -945 1305 -930
rect 1362 -945 1369 -930
rect 1479 -945 1486 -930
rect 1543 -945 1550 -930
rect 68 -1231 75 -1216
rect 132 -1231 139 -1216
rect 241 -1237 249 -1221
rect 351 -1235 358 -1220
rect 415 -1235 422 -1220
rect 611 -1215 617 -1204
rect 652 -1215 658 -1204
rect 703 -1215 709 -1204
rect 524 -1241 532 -1225
rect 196 -1563 203 -1548
rect 260 -1563 267 -1548
rect 399 -1563 406 -1548
rect 463 -1563 470 -1548
rect 586 -1563 595 -1548
rect 650 -1563 657 -1548
rect 767 -1563 774 -1548
rect 831 -1563 838 -1548
rect 936 -1569 943 -1554
rect 1000 -1569 1007 -1554
rect 1139 -1569 1146 -1554
rect 1203 -1569 1210 -1554
rect 1326 -1569 1333 -1554
rect 1390 -1569 1397 -1554
rect 1507 -1569 1514 -1554
rect 1571 -1569 1578 -1554
rect 96 -1855 103 -1840
rect 160 -1855 167 -1840
rect 269 -1861 277 -1845
rect 379 -1859 386 -1844
rect 443 -1859 450 -1844
rect 639 -1839 645 -1828
rect 680 -1839 686 -1828
rect 731 -1839 737 -1828
rect 552 -1865 560 -1849
<< ptransistor >>
rect -963 739 -956 754
rect -899 739 -892 754
rect -760 739 -753 754
rect -696 739 -689 754
rect -573 739 -566 754
rect -509 739 -502 754
rect -392 739 -385 754
rect -328 739 -321 754
rect -935 392 -928 407
rect -871 392 -864 407
rect -732 392 -725 407
rect -668 392 -661 407
rect -545 392 -538 407
rect -481 392 -474 407
rect -364 392 -357 407
rect -300 392 -293 407
rect -935 6 -928 21
rect -871 6 -864 21
rect -732 6 -725 21
rect -668 6 -661 21
rect -545 6 -538 21
rect -481 6 -474 21
rect -364 6 -357 21
rect -300 6 -293 21
rect -935 -418 -928 -403
rect -871 -418 -864 -403
rect -732 -418 -725 -403
rect -668 -418 -661 -403
rect -545 -418 -538 -403
rect -481 -418 -474 -403
rect -364 -418 -357 -403
rect -300 -418 -293 -403
rect 131 460 138 475
rect 195 460 202 475
rect 334 460 341 475
rect 398 460 405 475
rect 521 460 528 475
rect 585 460 592 475
rect 702 460 709 475
rect 766 460 773 475
rect 871 454 878 469
rect 935 454 942 469
rect 1074 454 1081 469
rect 1138 454 1145 469
rect 1261 454 1268 469
rect 1325 454 1332 469
rect 1442 454 1449 469
rect 1506 454 1513 469
rect 31 168 38 183
rect 95 168 103 183
rect 204 155 212 171
rect 314 164 321 179
rect 378 164 385 179
rect 487 151 495 167
rect 574 160 580 171
rect 615 160 621 171
rect 666 160 672 171
rect 188 -264 195 -249
rect 252 -264 259 -249
rect 391 -264 398 -249
rect 455 -264 462 -249
rect 578 -264 585 -249
rect 642 -264 649 -249
rect 759 -264 766 -249
rect 823 -264 830 -249
rect 928 -270 935 -255
rect 992 -270 999 -255
rect 1131 -270 1138 -255
rect 1195 -270 1202 -255
rect 1318 -270 1325 -255
rect 1382 -270 1389 -255
rect 1499 -270 1506 -255
rect 1563 -270 1570 -255
rect 88 -556 95 -541
rect 152 -556 160 -541
rect 261 -569 269 -553
rect 371 -560 378 -545
rect 435 -560 442 -545
rect 544 -573 552 -557
rect 631 -564 637 -553
rect 672 -564 678 -553
rect 723 -564 729 -553
rect 168 -854 175 -839
rect 232 -854 239 -839
rect 371 -854 378 -839
rect 435 -854 442 -839
rect 558 -854 565 -839
rect 622 -854 629 -839
rect 739 -854 746 -839
rect 803 -854 810 -839
rect 908 -860 915 -845
rect 972 -860 979 -845
rect 1111 -860 1118 -845
rect 1175 -860 1182 -845
rect 1298 -860 1305 -845
rect 1362 -860 1369 -845
rect 1479 -860 1486 -845
rect 1543 -860 1550 -845
rect 68 -1146 75 -1131
rect 132 -1146 140 -1131
rect 241 -1159 249 -1143
rect 351 -1150 358 -1135
rect 415 -1150 422 -1135
rect 524 -1163 532 -1147
rect 611 -1154 617 -1143
rect 652 -1154 658 -1143
rect 703 -1154 709 -1143
rect 196 -1478 203 -1463
rect 260 -1478 267 -1463
rect 399 -1478 406 -1463
rect 463 -1478 470 -1463
rect 586 -1478 593 -1463
rect 650 -1478 657 -1463
rect 767 -1478 774 -1463
rect 831 -1478 838 -1463
rect 936 -1484 943 -1469
rect 1000 -1484 1007 -1469
rect 1139 -1484 1146 -1469
rect 1203 -1484 1210 -1469
rect 1326 -1484 1333 -1469
rect 1390 -1484 1397 -1469
rect 1507 -1484 1514 -1469
rect 1571 -1484 1578 -1469
rect 96 -1770 103 -1755
rect 160 -1770 168 -1755
rect 269 -1783 277 -1767
rect 379 -1774 386 -1759
rect 443 -1774 450 -1759
rect 552 -1787 560 -1771
rect 639 -1778 645 -1767
rect 680 -1778 686 -1767
rect 731 -1778 737 -1767
<< ndiffusion >>
rect -977 667 -963 669
rect -977 660 -975 667
rect -967 660 -963 667
rect -977 654 -963 660
rect -956 666 -937 669
rect -956 657 -953 666
rect -943 657 -937 666
rect -956 654 -937 657
rect -918 668 -899 669
rect -918 660 -912 668
rect -904 660 -899 668
rect -918 654 -899 660
rect -892 667 -878 669
rect -892 659 -889 667
rect -881 659 -878 667
rect -892 654 -878 659
rect -774 667 -760 669
rect -774 660 -772 667
rect -764 660 -760 667
rect -774 654 -760 660
rect -753 666 -734 669
rect -753 657 -750 666
rect -740 657 -734 666
rect -753 654 -734 657
rect -715 668 -696 669
rect -715 660 -709 668
rect -701 660 -696 668
rect -715 654 -696 660
rect -689 667 -675 669
rect -689 659 -686 667
rect -678 659 -675 667
rect -689 654 -675 659
rect -587 667 -573 669
rect -587 660 -585 667
rect -577 660 -573 667
rect -587 654 -573 660
rect -566 666 -547 669
rect -566 657 -563 666
rect -553 657 -547 666
rect -566 654 -547 657
rect -528 668 -509 669
rect -528 660 -522 668
rect -514 660 -509 668
rect -528 654 -509 660
rect -502 667 -488 669
rect -502 659 -499 667
rect -491 659 -488 667
rect -502 654 -488 659
rect -406 667 -392 669
rect -406 660 -404 667
rect -396 660 -392 667
rect -406 654 -392 660
rect -385 666 -366 669
rect -385 657 -382 666
rect -372 657 -366 666
rect -385 654 -366 657
rect -347 668 -328 669
rect -347 660 -341 668
rect -333 660 -328 668
rect -347 654 -328 660
rect -321 667 -307 669
rect -321 659 -318 667
rect -310 659 -307 667
rect -321 654 -307 659
rect -949 320 -935 322
rect -949 313 -947 320
rect -939 313 -935 320
rect -949 307 -935 313
rect -928 319 -909 322
rect -928 310 -925 319
rect -915 310 -909 319
rect -928 307 -909 310
rect -890 321 -871 322
rect -890 313 -884 321
rect -876 313 -871 321
rect -890 307 -871 313
rect -864 320 -850 322
rect -864 312 -861 320
rect -853 312 -850 320
rect -864 307 -850 312
rect -746 320 -732 322
rect -746 313 -744 320
rect -736 313 -732 320
rect -746 307 -732 313
rect -725 319 -706 322
rect -725 310 -722 319
rect -712 310 -706 319
rect -725 307 -706 310
rect -687 321 -668 322
rect -687 313 -681 321
rect -673 313 -668 321
rect -687 307 -668 313
rect -661 320 -647 322
rect -661 312 -658 320
rect -650 312 -647 320
rect -661 307 -647 312
rect -559 320 -545 322
rect -559 313 -557 320
rect -549 313 -545 320
rect -559 307 -545 313
rect -538 319 -519 322
rect -538 310 -535 319
rect -525 310 -519 319
rect -538 307 -519 310
rect -500 321 -481 322
rect -500 313 -494 321
rect -486 313 -481 321
rect -500 307 -481 313
rect -474 320 -460 322
rect -474 312 -471 320
rect -463 312 -460 320
rect -474 307 -460 312
rect -378 320 -364 322
rect -378 313 -376 320
rect -368 313 -364 320
rect -378 307 -364 313
rect -357 319 -338 322
rect -357 310 -354 319
rect -344 310 -338 319
rect -357 307 -338 310
rect -319 321 -300 322
rect -319 313 -313 321
rect -305 313 -300 321
rect -319 307 -300 313
rect -293 320 -279 322
rect -293 312 -290 320
rect -282 312 -279 320
rect -293 307 -279 312
rect -949 -66 -935 -64
rect -949 -73 -947 -66
rect -939 -73 -935 -66
rect -949 -79 -935 -73
rect -928 -67 -909 -64
rect -928 -76 -925 -67
rect -915 -76 -909 -67
rect -928 -79 -909 -76
rect -890 -65 -871 -64
rect -890 -73 -884 -65
rect -876 -73 -871 -65
rect -890 -79 -871 -73
rect -864 -66 -850 -64
rect -864 -74 -861 -66
rect -853 -74 -850 -66
rect -864 -79 -850 -74
rect -746 -66 -732 -64
rect -746 -73 -744 -66
rect -736 -73 -732 -66
rect -746 -79 -732 -73
rect -725 -67 -706 -64
rect -725 -76 -722 -67
rect -712 -76 -706 -67
rect -725 -79 -706 -76
rect -687 -65 -668 -64
rect -687 -73 -681 -65
rect -673 -73 -668 -65
rect -687 -79 -668 -73
rect -661 -66 -647 -64
rect -661 -74 -658 -66
rect -650 -74 -647 -66
rect -661 -79 -647 -74
rect -559 -66 -545 -64
rect -559 -73 -557 -66
rect -549 -73 -545 -66
rect -559 -79 -545 -73
rect -538 -67 -519 -64
rect -538 -76 -535 -67
rect -525 -76 -519 -67
rect -538 -79 -519 -76
rect -500 -65 -481 -64
rect -500 -73 -494 -65
rect -486 -73 -481 -65
rect -500 -79 -481 -73
rect -474 -66 -460 -64
rect -474 -74 -471 -66
rect -463 -74 -460 -66
rect -474 -79 -460 -74
rect -378 -66 -364 -64
rect -378 -73 -376 -66
rect -368 -73 -364 -66
rect -378 -79 -364 -73
rect -357 -67 -338 -64
rect -357 -76 -354 -67
rect -344 -76 -338 -67
rect -357 -79 -338 -76
rect -319 -65 -300 -64
rect -319 -73 -313 -65
rect -305 -73 -300 -65
rect -319 -79 -300 -73
rect -293 -66 -279 -64
rect -293 -74 -290 -66
rect -282 -74 -279 -66
rect -293 -79 -279 -74
rect -949 -490 -935 -488
rect -949 -497 -947 -490
rect -939 -497 -935 -490
rect -949 -503 -935 -497
rect -928 -491 -909 -488
rect -928 -500 -925 -491
rect -915 -500 -909 -491
rect -928 -503 -909 -500
rect -890 -489 -871 -488
rect -890 -497 -884 -489
rect -876 -497 -871 -489
rect -890 -503 -871 -497
rect -864 -490 -850 -488
rect -864 -498 -861 -490
rect -853 -498 -850 -490
rect -864 -503 -850 -498
rect -746 -490 -732 -488
rect -746 -497 -744 -490
rect -736 -497 -732 -490
rect -746 -503 -732 -497
rect -725 -491 -706 -488
rect -725 -500 -722 -491
rect -712 -500 -706 -491
rect -725 -503 -706 -500
rect -687 -489 -668 -488
rect -687 -497 -681 -489
rect -673 -497 -668 -489
rect -687 -503 -668 -497
rect -661 -490 -647 -488
rect -661 -498 -658 -490
rect -650 -498 -647 -490
rect -661 -503 -647 -498
rect -559 -490 -545 -488
rect -559 -497 -557 -490
rect -549 -497 -545 -490
rect -559 -503 -545 -497
rect -538 -491 -519 -488
rect -538 -500 -535 -491
rect -525 -500 -519 -491
rect -538 -503 -519 -500
rect -500 -489 -481 -488
rect -500 -497 -494 -489
rect -486 -497 -481 -489
rect -500 -503 -481 -497
rect -474 -490 -460 -488
rect -474 -498 -471 -490
rect -463 -498 -460 -490
rect -474 -503 -460 -498
rect -378 -490 -364 -488
rect -378 -497 -376 -490
rect -368 -497 -364 -490
rect -378 -503 -364 -497
rect -357 -491 -338 -488
rect -357 -500 -354 -491
rect -344 -500 -338 -491
rect -357 -503 -338 -500
rect -319 -489 -300 -488
rect -319 -497 -313 -489
rect -305 -497 -300 -489
rect -319 -503 -300 -497
rect -293 -490 -279 -488
rect -293 -498 -290 -490
rect -282 -498 -279 -490
rect -293 -503 -279 -498
rect 117 388 131 390
rect 117 381 119 388
rect 127 381 131 388
rect 117 375 131 381
rect 138 387 157 390
rect 138 378 141 387
rect 151 378 157 387
rect 138 375 157 378
rect 176 389 195 390
rect 176 381 182 389
rect 190 381 195 389
rect 176 375 195 381
rect 202 388 216 390
rect 202 380 205 388
rect 213 380 216 388
rect 202 375 216 380
rect 320 388 334 390
rect 320 381 322 388
rect 330 381 334 388
rect 320 375 334 381
rect 341 387 360 390
rect 341 378 344 387
rect 354 378 360 387
rect 341 375 360 378
rect 379 389 398 390
rect 379 381 385 389
rect 393 381 398 389
rect 379 375 398 381
rect 405 388 419 390
rect 405 380 408 388
rect 416 380 419 388
rect 405 375 419 380
rect 507 388 521 390
rect 507 381 509 388
rect 517 381 521 388
rect 507 375 521 381
rect 530 387 547 390
rect 530 378 531 387
rect 541 378 547 387
rect 530 375 547 378
rect 566 389 585 390
rect 566 381 572 389
rect 580 381 585 389
rect 566 375 585 381
rect 592 388 606 390
rect 592 380 595 388
rect 603 380 606 388
rect 592 375 606 380
rect 688 388 702 390
rect 688 381 690 388
rect 698 381 702 388
rect 688 375 702 381
rect 709 387 728 390
rect 709 378 712 387
rect 722 378 728 387
rect 709 375 728 378
rect 747 389 766 390
rect 747 381 753 389
rect 761 381 766 389
rect 747 375 766 381
rect 773 388 787 390
rect 773 380 776 388
rect 784 380 787 388
rect 773 375 787 380
rect 857 382 871 384
rect 857 375 859 382
rect 867 375 871 382
rect 857 369 871 375
rect 878 381 897 384
rect 878 372 881 381
rect 891 372 897 381
rect 878 369 897 372
rect 916 383 935 384
rect 916 375 922 383
rect 930 375 935 383
rect 916 369 935 375
rect 942 382 956 384
rect 942 374 945 382
rect 953 374 956 382
rect 942 369 956 374
rect 1060 382 1074 384
rect 1060 375 1062 382
rect 1070 375 1074 382
rect 1060 369 1074 375
rect 1081 381 1100 384
rect 1081 372 1084 381
rect 1094 372 1100 381
rect 1081 369 1100 372
rect 1119 383 1138 384
rect 1119 375 1125 383
rect 1133 375 1138 383
rect 1119 369 1138 375
rect 1145 382 1159 384
rect 1145 374 1148 382
rect 1156 374 1159 382
rect 1145 369 1159 374
rect 1247 382 1261 384
rect 1247 375 1249 382
rect 1257 375 1261 382
rect 1247 369 1261 375
rect 1268 381 1287 384
rect 1268 372 1271 381
rect 1281 372 1287 381
rect 1268 369 1287 372
rect 1306 383 1325 384
rect 1306 375 1312 383
rect 1320 375 1325 383
rect 1306 369 1325 375
rect 1332 382 1346 384
rect 1332 374 1335 382
rect 1343 374 1346 382
rect 1332 369 1346 374
rect 1428 382 1442 384
rect 1428 375 1430 382
rect 1438 375 1442 382
rect 1428 369 1442 375
rect 1449 381 1468 384
rect 1449 372 1452 381
rect 1462 372 1468 381
rect 1449 369 1468 372
rect 1487 383 1506 384
rect 1487 375 1493 383
rect 1501 375 1506 383
rect 1487 369 1506 375
rect 1513 382 1527 384
rect 1513 374 1516 382
rect 1524 374 1527 382
rect 1513 369 1527 374
rect 17 96 31 98
rect 17 89 19 96
rect 27 89 31 96
rect 17 83 31 89
rect 38 95 57 98
rect 38 86 41 95
rect 51 86 57 95
rect 38 83 57 86
rect 76 97 95 98
rect 76 89 82 97
rect 90 89 95 97
rect 76 83 95 89
rect 102 96 116 98
rect 102 88 105 96
rect 113 88 116 96
rect 102 83 116 88
rect 187 89 204 93
rect 187 79 189 89
rect 199 79 204 89
rect 187 77 204 79
rect 212 90 227 93
rect 212 80 214 90
rect 224 80 227 90
rect 212 77 227 80
rect 300 92 314 94
rect 300 85 302 92
rect 310 85 314 92
rect 300 79 314 85
rect 321 91 340 94
rect 321 82 324 91
rect 334 82 340 91
rect 321 79 340 82
rect 359 93 378 94
rect 359 85 365 93
rect 373 85 378 93
rect 359 79 378 85
rect 385 92 399 94
rect 385 84 388 92
rect 396 84 399 92
rect 563 107 574 110
rect 563 102 565 107
rect 571 102 574 107
rect 563 99 574 102
rect 580 108 596 110
rect 580 102 584 108
rect 591 102 596 108
rect 580 99 596 102
rect 601 107 615 110
rect 601 102 605 107
rect 611 102 615 107
rect 601 99 615 102
rect 621 108 634 110
rect 621 102 624 108
rect 631 102 634 108
rect 621 99 634 102
rect 650 107 666 110
rect 650 102 656 107
rect 662 102 666 107
rect 650 99 666 102
rect 672 108 683 110
rect 672 102 674 108
rect 681 102 683 108
rect 672 99 683 102
rect 385 79 399 84
rect 470 85 487 89
rect 470 75 472 85
rect 482 75 487 85
rect 470 73 487 75
rect 495 86 510 89
rect 495 76 497 86
rect 507 76 510 86
rect 495 73 510 76
rect 174 -336 188 -334
rect 174 -343 176 -336
rect 184 -343 188 -336
rect 174 -349 188 -343
rect 195 -337 214 -334
rect 195 -346 198 -337
rect 208 -346 214 -337
rect 195 -349 214 -346
rect 233 -335 252 -334
rect 233 -343 239 -335
rect 247 -343 252 -335
rect 233 -349 252 -343
rect 259 -336 273 -334
rect 259 -344 262 -336
rect 270 -344 273 -336
rect 259 -349 273 -344
rect 377 -336 391 -334
rect 377 -343 379 -336
rect 387 -343 391 -336
rect 377 -349 391 -343
rect 398 -337 417 -334
rect 398 -346 401 -337
rect 411 -346 417 -337
rect 398 -349 417 -346
rect 436 -335 455 -334
rect 436 -343 442 -335
rect 450 -343 455 -335
rect 436 -349 455 -343
rect 462 -336 476 -334
rect 462 -344 465 -336
rect 473 -344 476 -336
rect 462 -349 476 -344
rect 564 -336 578 -334
rect 564 -343 566 -336
rect 574 -343 578 -336
rect 564 -349 578 -343
rect 587 -337 604 -334
rect 587 -346 588 -337
rect 598 -346 604 -337
rect 587 -349 604 -346
rect 623 -335 642 -334
rect 623 -343 629 -335
rect 637 -343 642 -335
rect 623 -349 642 -343
rect 649 -336 663 -334
rect 649 -344 652 -336
rect 660 -344 663 -336
rect 649 -349 663 -344
rect 745 -336 759 -334
rect 745 -343 747 -336
rect 755 -343 759 -336
rect 745 -349 759 -343
rect 766 -337 785 -334
rect 766 -346 769 -337
rect 779 -346 785 -337
rect 766 -349 785 -346
rect 804 -335 823 -334
rect 804 -343 810 -335
rect 818 -343 823 -335
rect 804 -349 823 -343
rect 830 -336 844 -334
rect 830 -344 833 -336
rect 841 -344 844 -336
rect 830 -349 844 -344
rect 914 -342 928 -340
rect 914 -349 916 -342
rect 924 -349 928 -342
rect 914 -355 928 -349
rect 935 -343 954 -340
rect 935 -352 938 -343
rect 948 -352 954 -343
rect 935 -355 954 -352
rect 973 -341 992 -340
rect 973 -349 979 -341
rect 987 -349 992 -341
rect 973 -355 992 -349
rect 999 -342 1013 -340
rect 999 -350 1002 -342
rect 1010 -350 1013 -342
rect 999 -355 1013 -350
rect 1117 -342 1131 -340
rect 1117 -349 1119 -342
rect 1127 -349 1131 -342
rect 1117 -355 1131 -349
rect 1138 -343 1157 -340
rect 1138 -352 1141 -343
rect 1151 -352 1157 -343
rect 1138 -355 1157 -352
rect 1176 -341 1195 -340
rect 1176 -349 1182 -341
rect 1190 -349 1195 -341
rect 1176 -355 1195 -349
rect 1202 -342 1216 -340
rect 1202 -350 1205 -342
rect 1213 -350 1216 -342
rect 1202 -355 1216 -350
rect 1304 -342 1318 -340
rect 1304 -349 1306 -342
rect 1314 -349 1318 -342
rect 1304 -355 1318 -349
rect 1325 -343 1344 -340
rect 1325 -352 1328 -343
rect 1338 -352 1344 -343
rect 1325 -355 1344 -352
rect 1363 -341 1382 -340
rect 1363 -349 1369 -341
rect 1377 -349 1382 -341
rect 1363 -355 1382 -349
rect 1389 -342 1403 -340
rect 1389 -350 1392 -342
rect 1400 -350 1403 -342
rect 1389 -355 1403 -350
rect 1485 -342 1499 -340
rect 1485 -349 1487 -342
rect 1495 -349 1499 -342
rect 1485 -355 1499 -349
rect 1506 -343 1525 -340
rect 1506 -352 1509 -343
rect 1519 -352 1525 -343
rect 1506 -355 1525 -352
rect 1544 -341 1563 -340
rect 1544 -349 1550 -341
rect 1558 -349 1563 -341
rect 1544 -355 1563 -349
rect 1570 -342 1584 -340
rect 1570 -350 1573 -342
rect 1581 -350 1584 -342
rect 1570 -355 1584 -350
rect 74 -628 88 -626
rect 74 -635 76 -628
rect 84 -635 88 -628
rect 74 -641 88 -635
rect 95 -629 114 -626
rect 95 -638 98 -629
rect 108 -638 114 -629
rect 95 -641 114 -638
rect 133 -627 152 -626
rect 133 -635 139 -627
rect 147 -635 152 -627
rect 133 -641 152 -635
rect 159 -628 173 -626
rect 159 -636 162 -628
rect 170 -636 173 -628
rect 159 -641 173 -636
rect 244 -635 261 -631
rect 244 -645 246 -635
rect 256 -645 261 -635
rect 244 -647 261 -645
rect 269 -634 284 -631
rect 269 -644 271 -634
rect 281 -644 284 -634
rect 269 -647 284 -644
rect 357 -632 371 -630
rect 357 -639 359 -632
rect 367 -639 371 -632
rect 357 -645 371 -639
rect 378 -633 397 -630
rect 378 -642 381 -633
rect 391 -642 397 -633
rect 378 -645 397 -642
rect 416 -631 435 -630
rect 416 -639 422 -631
rect 430 -639 435 -631
rect 416 -645 435 -639
rect 442 -632 456 -630
rect 442 -640 445 -632
rect 453 -640 456 -632
rect 620 -617 631 -614
rect 620 -622 622 -617
rect 628 -622 631 -617
rect 620 -625 631 -622
rect 637 -616 653 -614
rect 637 -622 641 -616
rect 648 -622 653 -616
rect 637 -625 653 -622
rect 658 -617 672 -614
rect 658 -622 662 -617
rect 668 -622 672 -617
rect 658 -625 672 -622
rect 678 -616 691 -614
rect 678 -622 681 -616
rect 688 -622 691 -616
rect 678 -625 691 -622
rect 707 -617 723 -614
rect 707 -622 713 -617
rect 719 -622 723 -617
rect 707 -625 723 -622
rect 729 -616 740 -614
rect 729 -622 731 -616
rect 738 -622 740 -616
rect 729 -625 740 -622
rect 442 -645 456 -640
rect 527 -639 544 -635
rect 527 -649 529 -639
rect 539 -649 544 -639
rect 527 -651 544 -649
rect 552 -638 567 -635
rect 552 -648 554 -638
rect 564 -648 567 -638
rect 552 -651 567 -648
rect 154 -926 168 -924
rect 154 -933 156 -926
rect 164 -933 168 -926
rect 154 -939 168 -933
rect 175 -927 194 -924
rect 175 -936 178 -927
rect 188 -936 194 -927
rect 175 -939 194 -936
rect 213 -925 232 -924
rect 213 -933 219 -925
rect 227 -933 232 -925
rect 213 -939 232 -933
rect 239 -926 253 -924
rect 239 -934 242 -926
rect 250 -934 253 -926
rect 239 -939 253 -934
rect 357 -926 371 -924
rect 357 -933 359 -926
rect 367 -933 371 -926
rect 357 -939 371 -933
rect 378 -927 397 -924
rect 378 -936 381 -927
rect 391 -936 397 -927
rect 378 -939 397 -936
rect 416 -925 435 -924
rect 416 -933 422 -925
rect 430 -933 435 -925
rect 416 -939 435 -933
rect 442 -926 456 -924
rect 442 -934 445 -926
rect 453 -934 456 -926
rect 442 -939 456 -934
rect 544 -926 558 -924
rect 544 -933 546 -926
rect 554 -933 558 -926
rect 544 -939 558 -933
rect 567 -927 584 -924
rect 567 -936 568 -927
rect 578 -936 584 -927
rect 567 -939 584 -936
rect 603 -925 622 -924
rect 603 -933 609 -925
rect 617 -933 622 -925
rect 603 -939 622 -933
rect 629 -926 643 -924
rect 629 -934 632 -926
rect 640 -934 643 -926
rect 629 -939 643 -934
rect 725 -926 739 -924
rect 725 -933 727 -926
rect 735 -933 739 -926
rect 725 -939 739 -933
rect 746 -927 765 -924
rect 746 -936 749 -927
rect 759 -936 765 -927
rect 746 -939 765 -936
rect 784 -925 803 -924
rect 784 -933 790 -925
rect 798 -933 803 -925
rect 784 -939 803 -933
rect 810 -926 824 -924
rect 810 -934 813 -926
rect 821 -934 824 -926
rect 810 -939 824 -934
rect 894 -932 908 -930
rect 894 -939 896 -932
rect 904 -939 908 -932
rect 894 -945 908 -939
rect 915 -933 934 -930
rect 915 -942 918 -933
rect 928 -942 934 -933
rect 915 -945 934 -942
rect 953 -931 972 -930
rect 953 -939 959 -931
rect 967 -939 972 -931
rect 953 -945 972 -939
rect 979 -932 993 -930
rect 979 -940 982 -932
rect 990 -940 993 -932
rect 979 -945 993 -940
rect 1097 -932 1111 -930
rect 1097 -939 1099 -932
rect 1107 -939 1111 -932
rect 1097 -945 1111 -939
rect 1118 -933 1137 -930
rect 1118 -942 1121 -933
rect 1131 -942 1137 -933
rect 1118 -945 1137 -942
rect 1156 -931 1175 -930
rect 1156 -939 1162 -931
rect 1170 -939 1175 -931
rect 1156 -945 1175 -939
rect 1182 -932 1196 -930
rect 1182 -940 1185 -932
rect 1193 -940 1196 -932
rect 1182 -945 1196 -940
rect 1284 -932 1298 -930
rect 1284 -939 1286 -932
rect 1294 -939 1298 -932
rect 1284 -945 1298 -939
rect 1305 -933 1324 -930
rect 1305 -942 1308 -933
rect 1318 -942 1324 -933
rect 1305 -945 1324 -942
rect 1343 -931 1362 -930
rect 1343 -939 1349 -931
rect 1357 -939 1362 -931
rect 1343 -945 1362 -939
rect 1369 -932 1383 -930
rect 1369 -940 1372 -932
rect 1380 -940 1383 -932
rect 1369 -945 1383 -940
rect 1465 -932 1479 -930
rect 1465 -939 1467 -932
rect 1475 -939 1479 -932
rect 1465 -945 1479 -939
rect 1486 -933 1505 -930
rect 1486 -942 1489 -933
rect 1499 -942 1505 -933
rect 1486 -945 1505 -942
rect 1524 -931 1543 -930
rect 1524 -939 1530 -931
rect 1538 -939 1543 -931
rect 1524 -945 1543 -939
rect 1550 -932 1564 -930
rect 1550 -940 1553 -932
rect 1561 -940 1564 -932
rect 1550 -945 1564 -940
rect 54 -1218 68 -1216
rect 54 -1225 56 -1218
rect 64 -1225 68 -1218
rect 54 -1231 68 -1225
rect 75 -1219 94 -1216
rect 75 -1228 78 -1219
rect 88 -1228 94 -1219
rect 75 -1231 94 -1228
rect 113 -1217 132 -1216
rect 113 -1225 119 -1217
rect 127 -1225 132 -1217
rect 113 -1231 132 -1225
rect 139 -1218 153 -1216
rect 139 -1226 142 -1218
rect 150 -1226 153 -1218
rect 139 -1231 153 -1226
rect 224 -1225 241 -1221
rect 224 -1235 226 -1225
rect 236 -1235 241 -1225
rect 224 -1237 241 -1235
rect 249 -1224 264 -1221
rect 249 -1234 251 -1224
rect 261 -1234 264 -1224
rect 249 -1237 264 -1234
rect 337 -1222 351 -1220
rect 337 -1229 339 -1222
rect 347 -1229 351 -1222
rect 337 -1235 351 -1229
rect 358 -1223 377 -1220
rect 358 -1232 361 -1223
rect 371 -1232 377 -1223
rect 358 -1235 377 -1232
rect 396 -1221 415 -1220
rect 396 -1229 402 -1221
rect 410 -1229 415 -1221
rect 396 -1235 415 -1229
rect 422 -1222 436 -1220
rect 422 -1230 425 -1222
rect 433 -1230 436 -1222
rect 600 -1207 611 -1204
rect 600 -1212 602 -1207
rect 608 -1212 611 -1207
rect 600 -1215 611 -1212
rect 617 -1206 633 -1204
rect 617 -1212 621 -1206
rect 628 -1212 633 -1206
rect 617 -1215 633 -1212
rect 638 -1207 652 -1204
rect 638 -1212 642 -1207
rect 648 -1212 652 -1207
rect 638 -1215 652 -1212
rect 658 -1206 671 -1204
rect 658 -1212 661 -1206
rect 668 -1212 671 -1206
rect 658 -1215 671 -1212
rect 687 -1207 703 -1204
rect 687 -1212 693 -1207
rect 699 -1212 703 -1207
rect 687 -1215 703 -1212
rect 709 -1206 720 -1204
rect 709 -1212 711 -1206
rect 718 -1212 720 -1206
rect 709 -1215 720 -1212
rect 422 -1235 436 -1230
rect 507 -1229 524 -1225
rect 507 -1239 509 -1229
rect 519 -1239 524 -1229
rect 507 -1241 524 -1239
rect 532 -1228 547 -1225
rect 532 -1238 534 -1228
rect 544 -1238 547 -1228
rect 532 -1241 547 -1238
rect 182 -1550 196 -1548
rect 182 -1557 184 -1550
rect 192 -1557 196 -1550
rect 182 -1563 196 -1557
rect 203 -1551 222 -1548
rect 203 -1560 206 -1551
rect 216 -1560 222 -1551
rect 203 -1563 222 -1560
rect 241 -1549 260 -1548
rect 241 -1557 247 -1549
rect 255 -1557 260 -1549
rect 241 -1563 260 -1557
rect 267 -1550 281 -1548
rect 267 -1558 270 -1550
rect 278 -1558 281 -1550
rect 267 -1563 281 -1558
rect 385 -1550 399 -1548
rect 385 -1557 387 -1550
rect 395 -1557 399 -1550
rect 385 -1563 399 -1557
rect 406 -1551 425 -1548
rect 406 -1560 409 -1551
rect 419 -1560 425 -1551
rect 406 -1563 425 -1560
rect 444 -1549 463 -1548
rect 444 -1557 450 -1549
rect 458 -1557 463 -1549
rect 444 -1563 463 -1557
rect 470 -1550 484 -1548
rect 470 -1558 473 -1550
rect 481 -1558 484 -1550
rect 470 -1563 484 -1558
rect 572 -1550 586 -1548
rect 572 -1557 574 -1550
rect 582 -1557 586 -1550
rect 572 -1563 586 -1557
rect 595 -1551 612 -1548
rect 595 -1560 596 -1551
rect 606 -1560 612 -1551
rect 595 -1563 612 -1560
rect 631 -1549 650 -1548
rect 631 -1557 637 -1549
rect 645 -1557 650 -1549
rect 631 -1563 650 -1557
rect 657 -1550 671 -1548
rect 657 -1558 660 -1550
rect 668 -1558 671 -1550
rect 657 -1563 671 -1558
rect 753 -1550 767 -1548
rect 753 -1557 755 -1550
rect 763 -1557 767 -1550
rect 753 -1563 767 -1557
rect 774 -1551 793 -1548
rect 774 -1560 777 -1551
rect 787 -1560 793 -1551
rect 774 -1563 793 -1560
rect 812 -1549 831 -1548
rect 812 -1557 818 -1549
rect 826 -1557 831 -1549
rect 812 -1563 831 -1557
rect 838 -1550 852 -1548
rect 838 -1558 841 -1550
rect 849 -1558 852 -1550
rect 838 -1563 852 -1558
rect 922 -1556 936 -1554
rect 922 -1563 924 -1556
rect 932 -1563 936 -1556
rect 922 -1569 936 -1563
rect 943 -1557 962 -1554
rect 943 -1566 946 -1557
rect 956 -1566 962 -1557
rect 943 -1569 962 -1566
rect 981 -1555 1000 -1554
rect 981 -1563 987 -1555
rect 995 -1563 1000 -1555
rect 981 -1569 1000 -1563
rect 1007 -1556 1021 -1554
rect 1007 -1564 1010 -1556
rect 1018 -1564 1021 -1556
rect 1007 -1569 1021 -1564
rect 1125 -1556 1139 -1554
rect 1125 -1563 1127 -1556
rect 1135 -1563 1139 -1556
rect 1125 -1569 1139 -1563
rect 1146 -1557 1165 -1554
rect 1146 -1566 1149 -1557
rect 1159 -1566 1165 -1557
rect 1146 -1569 1165 -1566
rect 1184 -1555 1203 -1554
rect 1184 -1563 1190 -1555
rect 1198 -1563 1203 -1555
rect 1184 -1569 1203 -1563
rect 1210 -1556 1224 -1554
rect 1210 -1564 1213 -1556
rect 1221 -1564 1224 -1556
rect 1210 -1569 1224 -1564
rect 1312 -1556 1326 -1554
rect 1312 -1563 1314 -1556
rect 1322 -1563 1326 -1556
rect 1312 -1569 1326 -1563
rect 1333 -1557 1352 -1554
rect 1333 -1566 1336 -1557
rect 1346 -1566 1352 -1557
rect 1333 -1569 1352 -1566
rect 1371 -1555 1390 -1554
rect 1371 -1563 1377 -1555
rect 1385 -1563 1390 -1555
rect 1371 -1569 1390 -1563
rect 1397 -1556 1411 -1554
rect 1397 -1564 1400 -1556
rect 1408 -1564 1411 -1556
rect 1397 -1569 1411 -1564
rect 1493 -1556 1507 -1554
rect 1493 -1563 1495 -1556
rect 1503 -1563 1507 -1556
rect 1493 -1569 1507 -1563
rect 1514 -1557 1533 -1554
rect 1514 -1566 1517 -1557
rect 1527 -1566 1533 -1557
rect 1514 -1569 1533 -1566
rect 1552 -1555 1571 -1554
rect 1552 -1563 1558 -1555
rect 1566 -1563 1571 -1555
rect 1552 -1569 1571 -1563
rect 1578 -1556 1592 -1554
rect 1578 -1564 1581 -1556
rect 1589 -1564 1592 -1556
rect 1578 -1569 1592 -1564
rect 82 -1842 96 -1840
rect 82 -1849 84 -1842
rect 92 -1849 96 -1842
rect 82 -1855 96 -1849
rect 103 -1843 122 -1840
rect 103 -1852 106 -1843
rect 116 -1852 122 -1843
rect 103 -1855 122 -1852
rect 141 -1841 160 -1840
rect 141 -1849 147 -1841
rect 155 -1849 160 -1841
rect 141 -1855 160 -1849
rect 167 -1842 181 -1840
rect 167 -1850 170 -1842
rect 178 -1850 181 -1842
rect 167 -1855 181 -1850
rect 252 -1849 269 -1845
rect 252 -1859 254 -1849
rect 264 -1859 269 -1849
rect 252 -1861 269 -1859
rect 277 -1848 292 -1845
rect 277 -1858 279 -1848
rect 289 -1858 292 -1848
rect 277 -1861 292 -1858
rect 365 -1846 379 -1844
rect 365 -1853 367 -1846
rect 375 -1853 379 -1846
rect 365 -1859 379 -1853
rect 386 -1847 405 -1844
rect 386 -1856 389 -1847
rect 399 -1856 405 -1847
rect 386 -1859 405 -1856
rect 424 -1845 443 -1844
rect 424 -1853 430 -1845
rect 438 -1853 443 -1845
rect 424 -1859 443 -1853
rect 450 -1846 464 -1844
rect 450 -1854 453 -1846
rect 461 -1854 464 -1846
rect 628 -1831 639 -1828
rect 628 -1836 630 -1831
rect 636 -1836 639 -1831
rect 628 -1839 639 -1836
rect 645 -1830 661 -1828
rect 645 -1836 649 -1830
rect 656 -1836 661 -1830
rect 645 -1839 661 -1836
rect 666 -1831 680 -1828
rect 666 -1836 670 -1831
rect 676 -1836 680 -1831
rect 666 -1839 680 -1836
rect 686 -1830 699 -1828
rect 686 -1836 689 -1830
rect 696 -1836 699 -1830
rect 686 -1839 699 -1836
rect 715 -1831 731 -1828
rect 715 -1836 721 -1831
rect 727 -1836 731 -1831
rect 715 -1839 731 -1836
rect 737 -1830 748 -1828
rect 737 -1836 739 -1830
rect 746 -1836 748 -1830
rect 737 -1839 748 -1836
rect 450 -1859 464 -1854
rect 535 -1853 552 -1849
rect 535 -1863 537 -1853
rect 547 -1863 552 -1853
rect 535 -1865 552 -1863
rect 560 -1852 575 -1849
rect 560 -1862 562 -1852
rect 572 -1862 575 -1852
rect 560 -1865 575 -1862
<< pdiffusion >>
rect -977 752 -963 754
rect -977 746 -974 752
rect -967 746 -963 752
rect -977 739 -963 746
rect -956 750 -937 754
rect -956 742 -952 750
rect -943 742 -937 750
rect -956 739 -937 742
rect -910 750 -899 754
rect -910 743 -908 750
rect -900 743 -899 750
rect -910 739 -899 743
rect -892 748 -870 754
rect -892 742 -889 748
rect -881 742 -870 748
rect -892 739 -870 742
rect -774 752 -760 754
rect -774 746 -771 752
rect -764 746 -760 752
rect -774 739 -760 746
rect -753 750 -734 754
rect -753 742 -749 750
rect -740 742 -734 750
rect -753 739 -734 742
rect -707 750 -696 754
rect -707 743 -705 750
rect -697 743 -696 750
rect -707 739 -696 743
rect -689 748 -667 754
rect -689 742 -686 748
rect -678 742 -667 748
rect -689 739 -667 742
rect -587 752 -573 754
rect -587 746 -584 752
rect -577 746 -573 752
rect -587 739 -573 746
rect -566 750 -547 754
rect -566 742 -562 750
rect -553 742 -547 750
rect -566 739 -547 742
rect -520 750 -509 754
rect -520 743 -518 750
rect -510 743 -509 750
rect -520 739 -509 743
rect -502 748 -480 754
rect -502 742 -499 748
rect -491 742 -480 748
rect -502 739 -480 742
rect -406 752 -392 754
rect -406 746 -403 752
rect -396 746 -392 752
rect -406 739 -392 746
rect -385 750 -366 754
rect -385 742 -381 750
rect -372 742 -366 750
rect -385 739 -366 742
rect -339 750 -328 754
rect -339 743 -337 750
rect -329 743 -328 750
rect -339 739 -328 743
rect -321 748 -299 754
rect -321 742 -318 748
rect -310 742 -299 748
rect -321 739 -299 742
rect -949 405 -935 407
rect -949 399 -946 405
rect -939 399 -935 405
rect -949 392 -935 399
rect -928 403 -909 407
rect -928 395 -924 403
rect -915 395 -909 403
rect -928 392 -909 395
rect -882 403 -871 407
rect -882 396 -880 403
rect -872 396 -871 403
rect -882 392 -871 396
rect -864 401 -842 407
rect -864 395 -861 401
rect -853 395 -842 401
rect -864 392 -842 395
rect -746 405 -732 407
rect -746 399 -743 405
rect -736 399 -732 405
rect -746 392 -732 399
rect -725 403 -706 407
rect -725 395 -721 403
rect -712 395 -706 403
rect -725 392 -706 395
rect -679 403 -668 407
rect -679 396 -677 403
rect -669 396 -668 403
rect -679 392 -668 396
rect -661 401 -639 407
rect -661 395 -658 401
rect -650 395 -639 401
rect -661 392 -639 395
rect -559 405 -545 407
rect -559 399 -556 405
rect -549 399 -545 405
rect -559 392 -545 399
rect -538 403 -519 407
rect -538 395 -534 403
rect -525 395 -519 403
rect -538 392 -519 395
rect -492 403 -481 407
rect -492 396 -490 403
rect -482 396 -481 403
rect -492 392 -481 396
rect -474 401 -452 407
rect -474 395 -471 401
rect -463 395 -452 401
rect -474 392 -452 395
rect -378 405 -364 407
rect -378 399 -375 405
rect -368 399 -364 405
rect -378 392 -364 399
rect -357 403 -338 407
rect -357 395 -353 403
rect -344 395 -338 403
rect -357 392 -338 395
rect -311 403 -300 407
rect -311 396 -309 403
rect -301 396 -300 403
rect -311 392 -300 396
rect -293 401 -271 407
rect -293 395 -290 401
rect -282 395 -271 401
rect -293 392 -271 395
rect -949 19 -935 21
rect -949 13 -946 19
rect -939 13 -935 19
rect -949 6 -935 13
rect -928 17 -909 21
rect -928 9 -924 17
rect -915 9 -909 17
rect -928 6 -909 9
rect -882 17 -871 21
rect -882 10 -880 17
rect -872 10 -871 17
rect -882 6 -871 10
rect -864 15 -842 21
rect -864 9 -861 15
rect -853 9 -842 15
rect -864 6 -842 9
rect -746 19 -732 21
rect -746 13 -743 19
rect -736 13 -732 19
rect -746 6 -732 13
rect -725 17 -706 21
rect -725 9 -721 17
rect -712 9 -706 17
rect -725 6 -706 9
rect -679 17 -668 21
rect -679 10 -677 17
rect -669 10 -668 17
rect -679 6 -668 10
rect -661 15 -639 21
rect -661 9 -658 15
rect -650 9 -639 15
rect -661 6 -639 9
rect -559 19 -545 21
rect -559 13 -556 19
rect -549 13 -545 19
rect -559 6 -545 13
rect -538 17 -519 21
rect -538 9 -534 17
rect -525 9 -519 17
rect -538 6 -519 9
rect -492 17 -481 21
rect -492 10 -490 17
rect -482 10 -481 17
rect -492 6 -481 10
rect -474 15 -452 21
rect -474 9 -471 15
rect -463 9 -452 15
rect -474 6 -452 9
rect -378 19 -364 21
rect -378 13 -375 19
rect -368 13 -364 19
rect -378 6 -364 13
rect -357 17 -338 21
rect -357 9 -353 17
rect -344 9 -338 17
rect -357 6 -338 9
rect -311 17 -300 21
rect -311 10 -309 17
rect -301 10 -300 17
rect -311 6 -300 10
rect -293 15 -271 21
rect -293 9 -290 15
rect -282 9 -271 15
rect -293 6 -271 9
rect -949 -405 -935 -403
rect -949 -411 -946 -405
rect -939 -411 -935 -405
rect -949 -418 -935 -411
rect -928 -407 -909 -403
rect -928 -415 -924 -407
rect -915 -415 -909 -407
rect -928 -418 -909 -415
rect -882 -407 -871 -403
rect -882 -414 -880 -407
rect -872 -414 -871 -407
rect -882 -418 -871 -414
rect -864 -409 -842 -403
rect -864 -415 -861 -409
rect -853 -415 -842 -409
rect -864 -418 -842 -415
rect -746 -405 -732 -403
rect -746 -411 -743 -405
rect -736 -411 -732 -405
rect -746 -418 -732 -411
rect -725 -407 -706 -403
rect -725 -415 -721 -407
rect -712 -415 -706 -407
rect -725 -418 -706 -415
rect -679 -407 -668 -403
rect -679 -414 -677 -407
rect -669 -414 -668 -407
rect -679 -418 -668 -414
rect -661 -409 -639 -403
rect -661 -415 -658 -409
rect -650 -415 -639 -409
rect -661 -418 -639 -415
rect -559 -405 -545 -403
rect -559 -411 -556 -405
rect -549 -411 -545 -405
rect -559 -418 -545 -411
rect -538 -407 -519 -403
rect -538 -415 -534 -407
rect -525 -415 -519 -407
rect -538 -418 -519 -415
rect -492 -407 -481 -403
rect -492 -414 -490 -407
rect -482 -414 -481 -407
rect -492 -418 -481 -414
rect -474 -409 -452 -403
rect -474 -415 -471 -409
rect -463 -415 -452 -409
rect -474 -418 -452 -415
rect -378 -405 -364 -403
rect -378 -411 -375 -405
rect -368 -411 -364 -405
rect -378 -418 -364 -411
rect -357 -407 -338 -403
rect -357 -415 -353 -407
rect -344 -415 -338 -407
rect -357 -418 -338 -415
rect -311 -407 -300 -403
rect -311 -414 -309 -407
rect -301 -414 -300 -407
rect -311 -418 -300 -414
rect -293 -409 -271 -403
rect -293 -415 -290 -409
rect -282 -415 -271 -409
rect -293 -418 -271 -415
rect 117 473 131 475
rect 117 467 120 473
rect 127 467 131 473
rect 117 460 131 467
rect 138 471 157 475
rect 138 463 142 471
rect 151 463 157 471
rect 138 460 157 463
rect 184 471 195 475
rect 184 464 186 471
rect 194 464 195 471
rect 184 460 195 464
rect 202 469 224 475
rect 202 463 205 469
rect 213 463 224 469
rect 202 460 224 463
rect 320 473 334 475
rect 320 467 323 473
rect 330 467 334 473
rect 320 460 334 467
rect 341 471 360 475
rect 341 463 345 471
rect 354 463 360 471
rect 341 460 360 463
rect 387 471 398 475
rect 387 464 389 471
rect 397 464 398 471
rect 387 460 398 464
rect 405 469 427 475
rect 405 463 408 469
rect 416 463 427 469
rect 405 460 427 463
rect 507 473 521 475
rect 507 467 510 473
rect 517 467 521 473
rect 507 460 521 467
rect 528 471 547 475
rect 528 463 532 471
rect 541 463 547 471
rect 528 460 547 463
rect 574 471 585 475
rect 574 464 576 471
rect 584 464 585 471
rect 574 460 585 464
rect 592 469 614 475
rect 592 463 595 469
rect 603 463 614 469
rect 592 460 614 463
rect 688 473 702 475
rect 688 467 691 473
rect 698 467 702 473
rect 688 460 702 467
rect 709 471 728 475
rect 709 463 713 471
rect 722 463 728 471
rect 709 460 728 463
rect 755 471 766 475
rect 755 464 757 471
rect 765 464 766 471
rect 755 460 766 464
rect 773 469 795 475
rect 773 463 776 469
rect 784 463 795 469
rect 773 460 795 463
rect 857 467 871 469
rect 857 461 860 467
rect 867 461 871 467
rect 857 454 871 461
rect 878 465 897 469
rect 878 457 882 465
rect 891 457 897 465
rect 878 454 897 457
rect 924 465 935 469
rect 924 458 926 465
rect 934 458 935 465
rect 924 454 935 458
rect 942 463 964 469
rect 942 457 945 463
rect 953 457 964 463
rect 942 454 964 457
rect 1060 467 1074 469
rect 1060 461 1063 467
rect 1070 461 1074 467
rect 1060 454 1074 461
rect 1081 465 1100 469
rect 1081 457 1085 465
rect 1094 457 1100 465
rect 1081 454 1100 457
rect 1127 465 1138 469
rect 1127 458 1129 465
rect 1137 458 1138 465
rect 1127 454 1138 458
rect 1145 463 1167 469
rect 1145 457 1148 463
rect 1156 457 1167 463
rect 1145 454 1167 457
rect 1247 467 1261 469
rect 1247 461 1250 467
rect 1257 461 1261 467
rect 1247 454 1261 461
rect 1268 465 1287 469
rect 1268 457 1272 465
rect 1281 457 1287 465
rect 1268 454 1287 457
rect 1314 465 1325 469
rect 1314 458 1316 465
rect 1324 458 1325 465
rect 1314 454 1325 458
rect 1332 463 1354 469
rect 1332 457 1335 463
rect 1343 457 1354 463
rect 1332 454 1354 457
rect 1428 467 1442 469
rect 1428 461 1431 467
rect 1438 461 1442 467
rect 1428 454 1442 461
rect 1449 465 1468 469
rect 1449 457 1453 465
rect 1462 457 1468 465
rect 1449 454 1468 457
rect 1495 465 1506 469
rect 1495 458 1497 465
rect 1505 458 1506 465
rect 1495 454 1506 458
rect 1513 463 1535 469
rect 1513 457 1516 463
rect 1524 457 1535 463
rect 1513 454 1535 457
rect 17 181 31 183
rect 17 175 20 181
rect 27 175 31 181
rect 17 168 31 175
rect 38 179 57 183
rect 38 171 42 179
rect 51 171 57 179
rect 38 168 57 171
rect 84 179 95 183
rect 84 172 86 179
rect 94 172 95 179
rect 84 168 95 172
rect 103 177 124 183
rect 103 171 105 177
rect 113 171 124 177
rect 103 168 124 171
rect 188 161 190 171
rect 200 161 204 171
rect 188 155 204 161
rect 212 168 228 171
rect 212 158 214 168
rect 224 158 228 168
rect 212 155 228 158
rect 300 177 314 179
rect 300 171 303 177
rect 310 171 314 177
rect 300 164 314 171
rect 321 175 340 179
rect 321 167 325 175
rect 334 167 340 175
rect 321 164 340 167
rect 367 175 378 179
rect 367 168 369 175
rect 377 168 378 175
rect 367 164 378 168
rect 385 173 407 179
rect 385 167 388 173
rect 396 167 407 173
rect 563 169 574 171
rect 385 164 407 167
rect 471 157 473 167
rect 483 157 487 167
rect 471 151 487 157
rect 495 164 511 167
rect 495 154 497 164
rect 507 154 511 164
rect 563 163 565 169
rect 571 163 574 169
rect 563 160 574 163
rect 580 166 596 171
rect 580 160 584 166
rect 590 160 596 166
rect 601 166 615 171
rect 601 160 605 166
rect 611 160 615 166
rect 621 166 634 171
rect 621 160 625 166
rect 631 160 634 166
rect 653 169 666 171
rect 653 163 656 169
rect 662 163 666 169
rect 653 160 666 163
rect 672 167 686 171
rect 672 161 674 167
rect 681 161 686 167
rect 672 160 686 161
rect 495 151 511 154
rect 174 -251 188 -249
rect 174 -257 177 -251
rect 184 -257 188 -251
rect 174 -264 188 -257
rect 195 -253 214 -249
rect 195 -261 199 -253
rect 208 -261 214 -253
rect 195 -264 214 -261
rect 241 -253 252 -249
rect 241 -260 243 -253
rect 251 -260 252 -253
rect 241 -264 252 -260
rect 259 -255 281 -249
rect 259 -261 262 -255
rect 270 -261 281 -255
rect 259 -264 281 -261
rect 377 -251 391 -249
rect 377 -257 380 -251
rect 387 -257 391 -251
rect 377 -264 391 -257
rect 398 -253 417 -249
rect 398 -261 402 -253
rect 411 -261 417 -253
rect 398 -264 417 -261
rect 444 -253 455 -249
rect 444 -260 446 -253
rect 454 -260 455 -253
rect 444 -264 455 -260
rect 462 -255 484 -249
rect 462 -261 465 -255
rect 473 -261 484 -255
rect 462 -264 484 -261
rect 564 -251 578 -249
rect 564 -257 567 -251
rect 574 -257 578 -251
rect 564 -264 578 -257
rect 585 -253 604 -249
rect 585 -261 589 -253
rect 598 -261 604 -253
rect 585 -264 604 -261
rect 631 -253 642 -249
rect 631 -260 633 -253
rect 641 -260 642 -253
rect 631 -264 642 -260
rect 649 -255 671 -249
rect 649 -261 652 -255
rect 660 -261 671 -255
rect 649 -264 671 -261
rect 745 -251 759 -249
rect 745 -257 748 -251
rect 755 -257 759 -251
rect 745 -264 759 -257
rect 766 -253 785 -249
rect 766 -261 770 -253
rect 779 -261 785 -253
rect 766 -264 785 -261
rect 812 -253 823 -249
rect 812 -260 814 -253
rect 822 -260 823 -253
rect 812 -264 823 -260
rect 830 -255 852 -249
rect 830 -261 833 -255
rect 841 -261 852 -255
rect 830 -264 852 -261
rect 914 -257 928 -255
rect 914 -263 917 -257
rect 924 -263 928 -257
rect 914 -270 928 -263
rect 935 -259 954 -255
rect 935 -267 939 -259
rect 948 -267 954 -259
rect 935 -270 954 -267
rect 981 -259 992 -255
rect 981 -266 983 -259
rect 991 -266 992 -259
rect 981 -270 992 -266
rect 999 -261 1021 -255
rect 999 -267 1002 -261
rect 1010 -267 1021 -261
rect 999 -270 1021 -267
rect 1117 -257 1131 -255
rect 1117 -263 1120 -257
rect 1127 -263 1131 -257
rect 1117 -270 1131 -263
rect 1138 -259 1157 -255
rect 1138 -267 1142 -259
rect 1151 -267 1157 -259
rect 1138 -270 1157 -267
rect 1184 -259 1195 -255
rect 1184 -266 1186 -259
rect 1194 -266 1195 -259
rect 1184 -270 1195 -266
rect 1202 -261 1224 -255
rect 1202 -267 1205 -261
rect 1213 -267 1224 -261
rect 1202 -270 1224 -267
rect 1304 -257 1318 -255
rect 1304 -263 1307 -257
rect 1314 -263 1318 -257
rect 1304 -270 1318 -263
rect 1325 -259 1344 -255
rect 1325 -267 1329 -259
rect 1338 -267 1344 -259
rect 1325 -270 1344 -267
rect 1371 -259 1382 -255
rect 1371 -266 1373 -259
rect 1381 -266 1382 -259
rect 1371 -270 1382 -266
rect 1389 -261 1411 -255
rect 1389 -267 1392 -261
rect 1400 -267 1411 -261
rect 1389 -270 1411 -267
rect 1485 -257 1499 -255
rect 1485 -263 1488 -257
rect 1495 -263 1499 -257
rect 1485 -270 1499 -263
rect 1506 -259 1525 -255
rect 1506 -267 1510 -259
rect 1519 -267 1525 -259
rect 1506 -270 1525 -267
rect 1552 -259 1563 -255
rect 1552 -266 1554 -259
rect 1562 -266 1563 -259
rect 1552 -270 1563 -266
rect 1570 -261 1592 -255
rect 1570 -267 1573 -261
rect 1581 -267 1592 -261
rect 1570 -270 1592 -267
rect 74 -543 88 -541
rect 74 -549 77 -543
rect 84 -549 88 -543
rect 74 -556 88 -549
rect 95 -545 114 -541
rect 95 -553 99 -545
rect 108 -553 114 -545
rect 95 -556 114 -553
rect 141 -545 152 -541
rect 141 -552 143 -545
rect 151 -552 152 -545
rect 141 -556 152 -552
rect 160 -547 181 -541
rect 160 -553 162 -547
rect 170 -553 181 -547
rect 160 -556 181 -553
rect 245 -563 247 -553
rect 257 -563 261 -553
rect 245 -569 261 -563
rect 269 -556 285 -553
rect 269 -566 271 -556
rect 281 -566 285 -556
rect 269 -569 285 -566
rect 357 -547 371 -545
rect 357 -553 360 -547
rect 367 -553 371 -547
rect 357 -560 371 -553
rect 378 -549 397 -545
rect 378 -557 382 -549
rect 391 -557 397 -549
rect 378 -560 397 -557
rect 424 -549 435 -545
rect 424 -556 426 -549
rect 434 -556 435 -549
rect 424 -560 435 -556
rect 442 -551 464 -545
rect 442 -557 445 -551
rect 453 -557 464 -551
rect 620 -555 631 -553
rect 442 -560 464 -557
rect 528 -567 530 -557
rect 540 -567 544 -557
rect 528 -573 544 -567
rect 552 -560 568 -557
rect 552 -570 554 -560
rect 564 -570 568 -560
rect 620 -561 622 -555
rect 628 -561 631 -555
rect 620 -564 631 -561
rect 637 -558 653 -553
rect 637 -564 641 -558
rect 647 -564 653 -558
rect 658 -558 672 -553
rect 658 -564 662 -558
rect 668 -564 672 -558
rect 678 -558 691 -553
rect 678 -564 682 -558
rect 688 -564 691 -558
rect 710 -555 723 -553
rect 710 -561 713 -555
rect 719 -561 723 -555
rect 710 -564 723 -561
rect 729 -557 743 -553
rect 729 -563 731 -557
rect 738 -563 743 -557
rect 729 -564 743 -563
rect 552 -573 568 -570
rect 154 -841 168 -839
rect 154 -847 157 -841
rect 164 -847 168 -841
rect 154 -854 168 -847
rect 175 -843 194 -839
rect 175 -851 179 -843
rect 188 -851 194 -843
rect 175 -854 194 -851
rect 221 -843 232 -839
rect 221 -850 223 -843
rect 231 -850 232 -843
rect 221 -854 232 -850
rect 239 -845 261 -839
rect 239 -851 242 -845
rect 250 -851 261 -845
rect 239 -854 261 -851
rect 357 -841 371 -839
rect 357 -847 360 -841
rect 367 -847 371 -841
rect 357 -854 371 -847
rect 378 -843 397 -839
rect 378 -851 382 -843
rect 391 -851 397 -843
rect 378 -854 397 -851
rect 424 -843 435 -839
rect 424 -850 426 -843
rect 434 -850 435 -843
rect 424 -854 435 -850
rect 442 -845 464 -839
rect 442 -851 445 -845
rect 453 -851 464 -845
rect 442 -854 464 -851
rect 544 -841 558 -839
rect 544 -847 547 -841
rect 554 -847 558 -841
rect 544 -854 558 -847
rect 565 -843 584 -839
rect 565 -851 569 -843
rect 578 -851 584 -843
rect 565 -854 584 -851
rect 611 -843 622 -839
rect 611 -850 613 -843
rect 621 -850 622 -843
rect 611 -854 622 -850
rect 629 -845 651 -839
rect 629 -851 632 -845
rect 640 -851 651 -845
rect 629 -854 651 -851
rect 725 -841 739 -839
rect 725 -847 728 -841
rect 735 -847 739 -841
rect 725 -854 739 -847
rect 746 -843 765 -839
rect 746 -851 750 -843
rect 759 -851 765 -843
rect 746 -854 765 -851
rect 792 -843 803 -839
rect 792 -850 794 -843
rect 802 -850 803 -843
rect 792 -854 803 -850
rect 810 -845 832 -839
rect 810 -851 813 -845
rect 821 -851 832 -845
rect 810 -854 832 -851
rect 894 -847 908 -845
rect 894 -853 897 -847
rect 904 -853 908 -847
rect 894 -860 908 -853
rect 915 -849 934 -845
rect 915 -857 919 -849
rect 928 -857 934 -849
rect 915 -860 934 -857
rect 961 -849 972 -845
rect 961 -856 963 -849
rect 971 -856 972 -849
rect 961 -860 972 -856
rect 979 -851 1001 -845
rect 979 -857 982 -851
rect 990 -857 1001 -851
rect 979 -860 1001 -857
rect 1097 -847 1111 -845
rect 1097 -853 1100 -847
rect 1107 -853 1111 -847
rect 1097 -860 1111 -853
rect 1118 -849 1137 -845
rect 1118 -857 1122 -849
rect 1131 -857 1137 -849
rect 1118 -860 1137 -857
rect 1164 -849 1175 -845
rect 1164 -856 1166 -849
rect 1174 -856 1175 -849
rect 1164 -860 1175 -856
rect 1182 -851 1204 -845
rect 1182 -857 1185 -851
rect 1193 -857 1204 -851
rect 1182 -860 1204 -857
rect 1284 -847 1298 -845
rect 1284 -853 1287 -847
rect 1294 -853 1298 -847
rect 1284 -860 1298 -853
rect 1305 -849 1324 -845
rect 1305 -857 1309 -849
rect 1318 -857 1324 -849
rect 1305 -860 1324 -857
rect 1351 -849 1362 -845
rect 1351 -856 1353 -849
rect 1361 -856 1362 -849
rect 1351 -860 1362 -856
rect 1369 -851 1391 -845
rect 1369 -857 1372 -851
rect 1380 -857 1391 -851
rect 1369 -860 1391 -857
rect 1465 -847 1479 -845
rect 1465 -853 1468 -847
rect 1475 -853 1479 -847
rect 1465 -860 1479 -853
rect 1486 -849 1505 -845
rect 1486 -857 1490 -849
rect 1499 -857 1505 -849
rect 1486 -860 1505 -857
rect 1532 -849 1543 -845
rect 1532 -856 1534 -849
rect 1542 -856 1543 -849
rect 1532 -860 1543 -856
rect 1550 -851 1572 -845
rect 1550 -857 1553 -851
rect 1561 -857 1572 -851
rect 1550 -860 1572 -857
rect 54 -1133 68 -1131
rect 54 -1139 57 -1133
rect 64 -1139 68 -1133
rect 54 -1146 68 -1139
rect 75 -1135 94 -1131
rect 75 -1143 79 -1135
rect 88 -1143 94 -1135
rect 75 -1146 94 -1143
rect 121 -1135 132 -1131
rect 121 -1142 123 -1135
rect 131 -1142 132 -1135
rect 121 -1146 132 -1142
rect 140 -1137 161 -1131
rect 140 -1143 142 -1137
rect 150 -1143 161 -1137
rect 140 -1146 161 -1143
rect 225 -1153 227 -1143
rect 237 -1153 241 -1143
rect 225 -1159 241 -1153
rect 249 -1146 265 -1143
rect 249 -1156 251 -1146
rect 261 -1156 265 -1146
rect 249 -1159 265 -1156
rect 337 -1137 351 -1135
rect 337 -1143 340 -1137
rect 347 -1143 351 -1137
rect 337 -1150 351 -1143
rect 358 -1139 377 -1135
rect 358 -1147 362 -1139
rect 371 -1147 377 -1139
rect 358 -1150 377 -1147
rect 404 -1139 415 -1135
rect 404 -1146 406 -1139
rect 414 -1146 415 -1139
rect 404 -1150 415 -1146
rect 422 -1141 444 -1135
rect 422 -1147 425 -1141
rect 433 -1147 444 -1141
rect 600 -1145 611 -1143
rect 422 -1150 444 -1147
rect 508 -1157 510 -1147
rect 520 -1157 524 -1147
rect 508 -1163 524 -1157
rect 532 -1150 548 -1147
rect 532 -1160 534 -1150
rect 544 -1160 548 -1150
rect 600 -1151 602 -1145
rect 608 -1151 611 -1145
rect 600 -1154 611 -1151
rect 617 -1148 633 -1143
rect 617 -1154 621 -1148
rect 627 -1154 633 -1148
rect 638 -1148 652 -1143
rect 638 -1154 642 -1148
rect 648 -1154 652 -1148
rect 658 -1148 671 -1143
rect 658 -1154 662 -1148
rect 668 -1154 671 -1148
rect 690 -1145 703 -1143
rect 690 -1151 693 -1145
rect 699 -1151 703 -1145
rect 690 -1154 703 -1151
rect 709 -1147 723 -1143
rect 709 -1153 711 -1147
rect 718 -1153 723 -1147
rect 709 -1154 723 -1153
rect 532 -1163 548 -1160
rect 182 -1465 196 -1463
rect 182 -1471 185 -1465
rect 192 -1471 196 -1465
rect 182 -1478 196 -1471
rect 203 -1467 222 -1463
rect 203 -1475 207 -1467
rect 216 -1475 222 -1467
rect 203 -1478 222 -1475
rect 249 -1467 260 -1463
rect 249 -1474 251 -1467
rect 259 -1474 260 -1467
rect 249 -1478 260 -1474
rect 267 -1469 289 -1463
rect 267 -1475 270 -1469
rect 278 -1475 289 -1469
rect 267 -1478 289 -1475
rect 385 -1465 399 -1463
rect 385 -1471 388 -1465
rect 395 -1471 399 -1465
rect 385 -1478 399 -1471
rect 406 -1467 425 -1463
rect 406 -1475 410 -1467
rect 419 -1475 425 -1467
rect 406 -1478 425 -1475
rect 452 -1467 463 -1463
rect 452 -1474 454 -1467
rect 462 -1474 463 -1467
rect 452 -1478 463 -1474
rect 470 -1469 492 -1463
rect 470 -1475 473 -1469
rect 481 -1475 492 -1469
rect 470 -1478 492 -1475
rect 572 -1465 586 -1463
rect 572 -1471 575 -1465
rect 582 -1471 586 -1465
rect 572 -1478 586 -1471
rect 593 -1467 612 -1463
rect 593 -1475 597 -1467
rect 606 -1475 612 -1467
rect 593 -1478 612 -1475
rect 639 -1467 650 -1463
rect 639 -1474 641 -1467
rect 649 -1474 650 -1467
rect 639 -1478 650 -1474
rect 657 -1469 679 -1463
rect 657 -1475 660 -1469
rect 668 -1475 679 -1469
rect 657 -1478 679 -1475
rect 753 -1465 767 -1463
rect 753 -1471 756 -1465
rect 763 -1471 767 -1465
rect 753 -1478 767 -1471
rect 774 -1467 793 -1463
rect 774 -1475 778 -1467
rect 787 -1475 793 -1467
rect 774 -1478 793 -1475
rect 820 -1467 831 -1463
rect 820 -1474 822 -1467
rect 830 -1474 831 -1467
rect 820 -1478 831 -1474
rect 838 -1469 860 -1463
rect 838 -1475 841 -1469
rect 849 -1475 860 -1469
rect 838 -1478 860 -1475
rect 922 -1471 936 -1469
rect 922 -1477 925 -1471
rect 932 -1477 936 -1471
rect 922 -1484 936 -1477
rect 943 -1473 962 -1469
rect 943 -1481 947 -1473
rect 956 -1481 962 -1473
rect 943 -1484 962 -1481
rect 989 -1473 1000 -1469
rect 989 -1480 991 -1473
rect 999 -1480 1000 -1473
rect 989 -1484 1000 -1480
rect 1007 -1475 1029 -1469
rect 1007 -1481 1010 -1475
rect 1018 -1481 1029 -1475
rect 1007 -1484 1029 -1481
rect 1125 -1471 1139 -1469
rect 1125 -1477 1128 -1471
rect 1135 -1477 1139 -1471
rect 1125 -1484 1139 -1477
rect 1146 -1473 1165 -1469
rect 1146 -1481 1150 -1473
rect 1159 -1481 1165 -1473
rect 1146 -1484 1165 -1481
rect 1192 -1473 1203 -1469
rect 1192 -1480 1194 -1473
rect 1202 -1480 1203 -1473
rect 1192 -1484 1203 -1480
rect 1210 -1475 1232 -1469
rect 1210 -1481 1213 -1475
rect 1221 -1481 1232 -1475
rect 1210 -1484 1232 -1481
rect 1312 -1471 1326 -1469
rect 1312 -1477 1315 -1471
rect 1322 -1477 1326 -1471
rect 1312 -1484 1326 -1477
rect 1333 -1473 1352 -1469
rect 1333 -1481 1337 -1473
rect 1346 -1481 1352 -1473
rect 1333 -1484 1352 -1481
rect 1379 -1473 1390 -1469
rect 1379 -1480 1381 -1473
rect 1389 -1480 1390 -1473
rect 1379 -1484 1390 -1480
rect 1397 -1475 1419 -1469
rect 1397 -1481 1400 -1475
rect 1408 -1481 1419 -1475
rect 1397 -1484 1419 -1481
rect 1493 -1471 1507 -1469
rect 1493 -1477 1496 -1471
rect 1503 -1477 1507 -1471
rect 1493 -1484 1507 -1477
rect 1514 -1473 1533 -1469
rect 1514 -1481 1518 -1473
rect 1527 -1481 1533 -1473
rect 1514 -1484 1533 -1481
rect 1560 -1473 1571 -1469
rect 1560 -1480 1562 -1473
rect 1570 -1480 1571 -1473
rect 1560 -1484 1571 -1480
rect 1578 -1475 1600 -1469
rect 1578 -1481 1581 -1475
rect 1589 -1481 1600 -1475
rect 1578 -1484 1600 -1481
rect 82 -1757 96 -1755
rect 82 -1763 85 -1757
rect 92 -1763 96 -1757
rect 82 -1770 96 -1763
rect 103 -1759 122 -1755
rect 103 -1767 107 -1759
rect 116 -1767 122 -1759
rect 103 -1770 122 -1767
rect 149 -1759 160 -1755
rect 149 -1766 151 -1759
rect 159 -1766 160 -1759
rect 149 -1770 160 -1766
rect 168 -1761 189 -1755
rect 168 -1767 170 -1761
rect 178 -1767 189 -1761
rect 168 -1770 189 -1767
rect 253 -1777 255 -1767
rect 265 -1777 269 -1767
rect 253 -1783 269 -1777
rect 277 -1770 293 -1767
rect 277 -1780 279 -1770
rect 289 -1780 293 -1770
rect 277 -1783 293 -1780
rect 365 -1761 379 -1759
rect 365 -1767 368 -1761
rect 375 -1767 379 -1761
rect 365 -1774 379 -1767
rect 386 -1763 405 -1759
rect 386 -1771 390 -1763
rect 399 -1771 405 -1763
rect 386 -1774 405 -1771
rect 432 -1763 443 -1759
rect 432 -1770 434 -1763
rect 442 -1770 443 -1763
rect 432 -1774 443 -1770
rect 450 -1765 472 -1759
rect 450 -1771 453 -1765
rect 461 -1771 472 -1765
rect 628 -1769 639 -1767
rect 450 -1774 472 -1771
rect 536 -1781 538 -1771
rect 548 -1781 552 -1771
rect 536 -1787 552 -1781
rect 560 -1774 576 -1771
rect 560 -1784 562 -1774
rect 572 -1784 576 -1774
rect 628 -1775 630 -1769
rect 636 -1775 639 -1769
rect 628 -1778 639 -1775
rect 645 -1772 661 -1767
rect 645 -1778 649 -1772
rect 655 -1778 661 -1772
rect 666 -1772 680 -1767
rect 666 -1778 670 -1772
rect 676 -1778 680 -1772
rect 686 -1772 699 -1767
rect 686 -1778 690 -1772
rect 696 -1778 699 -1772
rect 718 -1769 731 -1767
rect 718 -1775 721 -1769
rect 727 -1775 731 -1769
rect 718 -1778 731 -1775
rect 737 -1771 751 -1767
rect 737 -1777 739 -1771
rect 746 -1777 751 -1771
rect 737 -1778 751 -1777
rect 560 -1787 576 -1784
<< ndcontact >>
rect -975 660 -967 667
rect -953 657 -943 666
rect -912 660 -904 668
rect -889 659 -881 667
rect -772 660 -764 667
rect -750 657 -740 666
rect -709 660 -701 668
rect -686 659 -678 667
rect -585 660 -577 667
rect -563 657 -553 666
rect -522 660 -514 668
rect -499 659 -491 667
rect -404 660 -396 667
rect -382 657 -372 666
rect -341 660 -333 668
rect -318 659 -310 667
rect -947 313 -939 320
rect -925 310 -915 319
rect -884 313 -876 321
rect -861 312 -853 320
rect -744 313 -736 320
rect -722 310 -712 319
rect -681 313 -673 321
rect -658 312 -650 320
rect -557 313 -549 320
rect -535 310 -525 319
rect -494 313 -486 321
rect -471 312 -463 320
rect -376 313 -368 320
rect -354 310 -344 319
rect -313 313 -305 321
rect -290 312 -282 320
rect -947 -73 -939 -66
rect -925 -76 -915 -67
rect -884 -73 -876 -65
rect -861 -74 -853 -66
rect -744 -73 -736 -66
rect -722 -76 -712 -67
rect -681 -73 -673 -65
rect -658 -74 -650 -66
rect -557 -73 -549 -66
rect -535 -76 -525 -67
rect -494 -73 -486 -65
rect -471 -74 -463 -66
rect -376 -73 -368 -66
rect -354 -76 -344 -67
rect -313 -73 -305 -65
rect -290 -74 -282 -66
rect -947 -497 -939 -490
rect -925 -500 -915 -491
rect -884 -497 -876 -489
rect -861 -498 -853 -490
rect -744 -497 -736 -490
rect -722 -500 -712 -491
rect -681 -497 -673 -489
rect -658 -498 -650 -490
rect -557 -497 -549 -490
rect -535 -500 -525 -491
rect -494 -497 -486 -489
rect -471 -498 -463 -490
rect -376 -497 -368 -490
rect -354 -500 -344 -491
rect -313 -497 -305 -489
rect -290 -498 -282 -490
rect 119 381 127 388
rect 141 378 151 387
rect 182 381 190 389
rect 205 380 213 388
rect 322 381 330 388
rect 344 378 354 387
rect 385 381 393 389
rect 408 380 416 388
rect 509 381 517 388
rect 531 378 541 387
rect 572 381 580 389
rect 595 380 603 388
rect 690 381 698 388
rect 712 378 722 387
rect 753 381 761 389
rect 776 380 784 388
rect 859 375 867 382
rect 881 372 891 381
rect 922 375 930 383
rect 945 374 953 382
rect 1062 375 1070 382
rect 1084 372 1094 381
rect 1125 375 1133 383
rect 1148 374 1156 382
rect 1249 375 1257 382
rect 1271 372 1281 381
rect 1312 375 1320 383
rect 1335 374 1343 382
rect 1430 375 1438 382
rect 1452 372 1462 381
rect 1493 375 1501 383
rect 1516 374 1524 382
rect 19 89 27 96
rect 41 86 51 95
rect 82 89 90 97
rect 105 88 113 96
rect 189 79 199 89
rect 214 80 224 90
rect 302 85 310 92
rect 324 82 334 91
rect 365 85 373 93
rect 388 84 396 92
rect 565 102 571 107
rect 584 102 591 108
rect 605 102 611 107
rect 624 102 631 108
rect 656 102 662 107
rect 674 102 681 108
rect 472 75 482 85
rect 497 76 507 86
rect 176 -343 184 -336
rect 198 -346 208 -337
rect 239 -343 247 -335
rect 262 -344 270 -336
rect 379 -343 387 -336
rect 401 -346 411 -337
rect 442 -343 450 -335
rect 465 -344 473 -336
rect 566 -343 574 -336
rect 588 -346 598 -337
rect 629 -343 637 -335
rect 652 -344 660 -336
rect 747 -343 755 -336
rect 769 -346 779 -337
rect 810 -343 818 -335
rect 833 -344 841 -336
rect 916 -349 924 -342
rect 938 -352 948 -343
rect 979 -349 987 -341
rect 1002 -350 1010 -342
rect 1119 -349 1127 -342
rect 1141 -352 1151 -343
rect 1182 -349 1190 -341
rect 1205 -350 1213 -342
rect 1306 -349 1314 -342
rect 1328 -352 1338 -343
rect 1369 -349 1377 -341
rect 1392 -350 1400 -342
rect 1487 -349 1495 -342
rect 1509 -352 1519 -343
rect 1550 -349 1558 -341
rect 1573 -350 1581 -342
rect 76 -635 84 -628
rect 98 -638 108 -629
rect 139 -635 147 -627
rect 162 -636 170 -628
rect 246 -645 256 -635
rect 271 -644 281 -634
rect 359 -639 367 -632
rect 381 -642 391 -633
rect 422 -639 430 -631
rect 445 -640 453 -632
rect 622 -622 628 -617
rect 641 -622 648 -616
rect 662 -622 668 -617
rect 681 -622 688 -616
rect 713 -622 719 -617
rect 731 -622 738 -616
rect 529 -649 539 -639
rect 554 -648 564 -638
rect 156 -933 164 -926
rect 178 -936 188 -927
rect 219 -933 227 -925
rect 242 -934 250 -926
rect 359 -933 367 -926
rect 381 -936 391 -927
rect 422 -933 430 -925
rect 445 -934 453 -926
rect 546 -933 554 -926
rect 568 -936 578 -927
rect 609 -933 617 -925
rect 632 -934 640 -926
rect 727 -933 735 -926
rect 749 -936 759 -927
rect 790 -933 798 -925
rect 813 -934 821 -926
rect 896 -939 904 -932
rect 918 -942 928 -933
rect 959 -939 967 -931
rect 982 -940 990 -932
rect 1099 -939 1107 -932
rect 1121 -942 1131 -933
rect 1162 -939 1170 -931
rect 1185 -940 1193 -932
rect 1286 -939 1294 -932
rect 1308 -942 1318 -933
rect 1349 -939 1357 -931
rect 1372 -940 1380 -932
rect 1467 -939 1475 -932
rect 1489 -942 1499 -933
rect 1530 -939 1538 -931
rect 1553 -940 1561 -932
rect 56 -1225 64 -1218
rect 78 -1228 88 -1219
rect 119 -1225 127 -1217
rect 142 -1226 150 -1218
rect 226 -1235 236 -1225
rect 251 -1234 261 -1224
rect 339 -1229 347 -1222
rect 361 -1232 371 -1223
rect 402 -1229 410 -1221
rect 425 -1230 433 -1222
rect 602 -1212 608 -1207
rect 621 -1212 628 -1206
rect 642 -1212 648 -1207
rect 661 -1212 668 -1206
rect 693 -1212 699 -1207
rect 711 -1212 718 -1206
rect 509 -1239 519 -1229
rect 534 -1238 544 -1228
rect 184 -1557 192 -1550
rect 206 -1560 216 -1551
rect 247 -1557 255 -1549
rect 270 -1558 278 -1550
rect 387 -1557 395 -1550
rect 409 -1560 419 -1551
rect 450 -1557 458 -1549
rect 473 -1558 481 -1550
rect 574 -1557 582 -1550
rect 596 -1560 606 -1551
rect 637 -1557 645 -1549
rect 660 -1558 668 -1550
rect 755 -1557 763 -1550
rect 777 -1560 787 -1551
rect 818 -1557 826 -1549
rect 841 -1558 849 -1550
rect 924 -1563 932 -1556
rect 946 -1566 956 -1557
rect 987 -1563 995 -1555
rect 1010 -1564 1018 -1556
rect 1127 -1563 1135 -1556
rect 1149 -1566 1159 -1557
rect 1190 -1563 1198 -1555
rect 1213 -1564 1221 -1556
rect 1314 -1563 1322 -1556
rect 1336 -1566 1346 -1557
rect 1377 -1563 1385 -1555
rect 1400 -1564 1408 -1556
rect 1495 -1563 1503 -1556
rect 1517 -1566 1527 -1557
rect 1558 -1563 1566 -1555
rect 1581 -1564 1589 -1556
rect 84 -1849 92 -1842
rect 106 -1852 116 -1843
rect 147 -1849 155 -1841
rect 170 -1850 178 -1842
rect 254 -1859 264 -1849
rect 279 -1858 289 -1848
rect 367 -1853 375 -1846
rect 389 -1856 399 -1847
rect 430 -1853 438 -1845
rect 453 -1854 461 -1846
rect 630 -1836 636 -1831
rect 649 -1836 656 -1830
rect 670 -1836 676 -1831
rect 689 -1836 696 -1830
rect 721 -1836 727 -1831
rect 739 -1836 746 -1830
rect 537 -1863 547 -1853
rect 562 -1862 572 -1852
<< pdcontact >>
rect -974 746 -967 752
rect -952 742 -943 750
rect -908 743 -900 750
rect -889 742 -881 748
rect -771 746 -764 752
rect -749 742 -740 750
rect -705 743 -697 750
rect -686 742 -678 748
rect -584 746 -577 752
rect -562 742 -553 750
rect -518 743 -510 750
rect -499 742 -491 748
rect -403 746 -396 752
rect -381 742 -372 750
rect -337 743 -329 750
rect -318 742 -310 748
rect -946 399 -939 405
rect -924 395 -915 403
rect -880 396 -872 403
rect -861 395 -853 401
rect -743 399 -736 405
rect -721 395 -712 403
rect -677 396 -669 403
rect -658 395 -650 401
rect -556 399 -549 405
rect -534 395 -525 403
rect -490 396 -482 403
rect -471 395 -463 401
rect -375 399 -368 405
rect -353 395 -344 403
rect -309 396 -301 403
rect -290 395 -282 401
rect -946 13 -939 19
rect -924 9 -915 17
rect -880 10 -872 17
rect -861 9 -853 15
rect -743 13 -736 19
rect -721 9 -712 17
rect -677 10 -669 17
rect -658 9 -650 15
rect -556 13 -549 19
rect -534 9 -525 17
rect -490 10 -482 17
rect -471 9 -463 15
rect -375 13 -368 19
rect -353 9 -344 17
rect -309 10 -301 17
rect -290 9 -282 15
rect -946 -411 -939 -405
rect -924 -415 -915 -407
rect -880 -414 -872 -407
rect -861 -415 -853 -409
rect -743 -411 -736 -405
rect -721 -415 -712 -407
rect -677 -414 -669 -407
rect -658 -415 -650 -409
rect -556 -411 -549 -405
rect -534 -415 -525 -407
rect -490 -414 -482 -407
rect -471 -415 -463 -409
rect -375 -411 -368 -405
rect -353 -415 -344 -407
rect -309 -414 -301 -407
rect -290 -415 -282 -409
rect 120 467 127 473
rect 142 463 151 471
rect 186 464 194 471
rect 205 463 213 469
rect 323 467 330 473
rect 345 463 354 471
rect 389 464 397 471
rect 408 463 416 469
rect 510 467 517 473
rect 532 463 541 471
rect 576 464 584 471
rect 595 463 603 469
rect 691 467 698 473
rect 713 463 722 471
rect 757 464 765 471
rect 776 463 784 469
rect 860 461 867 467
rect 882 457 891 465
rect 926 458 934 465
rect 945 457 953 463
rect 1063 461 1070 467
rect 1085 457 1094 465
rect 1129 458 1137 465
rect 1148 457 1156 463
rect 1250 461 1257 467
rect 1272 457 1281 465
rect 1316 458 1324 465
rect 1335 457 1343 463
rect 1431 461 1438 467
rect 1453 457 1462 465
rect 1497 458 1505 465
rect 1516 457 1524 463
rect 20 175 27 181
rect 42 171 51 179
rect 86 172 94 179
rect 105 171 113 177
rect 190 161 200 171
rect 214 158 224 168
rect 303 171 310 177
rect 325 167 334 175
rect 369 168 377 175
rect 388 167 396 173
rect 473 157 483 167
rect 497 154 507 164
rect 565 163 571 169
rect 584 160 590 166
rect 605 160 611 166
rect 625 160 631 166
rect 656 163 662 169
rect 674 161 681 167
rect 177 -257 184 -251
rect 199 -261 208 -253
rect 243 -260 251 -253
rect 262 -261 270 -255
rect 380 -257 387 -251
rect 402 -261 411 -253
rect 446 -260 454 -253
rect 465 -261 473 -255
rect 567 -257 574 -251
rect 589 -261 598 -253
rect 633 -260 641 -253
rect 652 -261 660 -255
rect 748 -257 755 -251
rect 770 -261 779 -253
rect 814 -260 822 -253
rect 833 -261 841 -255
rect 917 -263 924 -257
rect 939 -267 948 -259
rect 983 -266 991 -259
rect 1002 -267 1010 -261
rect 1120 -263 1127 -257
rect 1142 -267 1151 -259
rect 1186 -266 1194 -259
rect 1205 -267 1213 -261
rect 1307 -263 1314 -257
rect 1329 -267 1338 -259
rect 1373 -266 1381 -259
rect 1392 -267 1400 -261
rect 1488 -263 1495 -257
rect 1510 -267 1519 -259
rect 1554 -266 1562 -259
rect 1573 -267 1581 -261
rect 77 -549 84 -543
rect 99 -553 108 -545
rect 143 -552 151 -545
rect 162 -553 170 -547
rect 247 -563 257 -553
rect 271 -566 281 -556
rect 360 -553 367 -547
rect 382 -557 391 -549
rect 426 -556 434 -549
rect 445 -557 453 -551
rect 530 -567 540 -557
rect 554 -570 564 -560
rect 622 -561 628 -555
rect 641 -564 647 -558
rect 662 -564 668 -558
rect 682 -564 688 -558
rect 713 -561 719 -555
rect 731 -563 738 -557
rect 157 -847 164 -841
rect 179 -851 188 -843
rect 223 -850 231 -843
rect 242 -851 250 -845
rect 360 -847 367 -841
rect 382 -851 391 -843
rect 426 -850 434 -843
rect 445 -851 453 -845
rect 547 -847 554 -841
rect 569 -851 578 -843
rect 613 -850 621 -843
rect 632 -851 640 -845
rect 728 -847 735 -841
rect 750 -851 759 -843
rect 794 -850 802 -843
rect 813 -851 821 -845
rect 897 -853 904 -847
rect 919 -857 928 -849
rect 963 -856 971 -849
rect 982 -857 990 -851
rect 1100 -853 1107 -847
rect 1122 -857 1131 -849
rect 1166 -856 1174 -849
rect 1185 -857 1193 -851
rect 1287 -853 1294 -847
rect 1309 -857 1318 -849
rect 1353 -856 1361 -849
rect 1372 -857 1380 -851
rect 1468 -853 1475 -847
rect 1490 -857 1499 -849
rect 1534 -856 1542 -849
rect 1553 -857 1561 -851
rect 57 -1139 64 -1133
rect 79 -1143 88 -1135
rect 123 -1142 131 -1135
rect 142 -1143 150 -1137
rect 227 -1153 237 -1143
rect 251 -1156 261 -1146
rect 340 -1143 347 -1137
rect 362 -1147 371 -1139
rect 406 -1146 414 -1139
rect 425 -1147 433 -1141
rect 510 -1157 520 -1147
rect 534 -1160 544 -1150
rect 602 -1151 608 -1145
rect 621 -1154 627 -1148
rect 642 -1154 648 -1148
rect 662 -1154 668 -1148
rect 693 -1151 699 -1145
rect 711 -1153 718 -1147
rect 185 -1471 192 -1465
rect 207 -1475 216 -1467
rect 251 -1474 259 -1467
rect 270 -1475 278 -1469
rect 388 -1471 395 -1465
rect 410 -1475 419 -1467
rect 454 -1474 462 -1467
rect 473 -1475 481 -1469
rect 575 -1471 582 -1465
rect 597 -1475 606 -1467
rect 641 -1474 649 -1467
rect 660 -1475 668 -1469
rect 756 -1471 763 -1465
rect 778 -1475 787 -1467
rect 822 -1474 830 -1467
rect 841 -1475 849 -1469
rect 925 -1477 932 -1471
rect 947 -1481 956 -1473
rect 991 -1480 999 -1473
rect 1010 -1481 1018 -1475
rect 1128 -1477 1135 -1471
rect 1150 -1481 1159 -1473
rect 1194 -1480 1202 -1473
rect 1213 -1481 1221 -1475
rect 1315 -1477 1322 -1471
rect 1337 -1481 1346 -1473
rect 1381 -1480 1389 -1473
rect 1400 -1481 1408 -1475
rect 1496 -1477 1503 -1471
rect 1518 -1481 1527 -1473
rect 1562 -1480 1570 -1473
rect 1581 -1481 1589 -1475
rect 85 -1763 92 -1757
rect 107 -1767 116 -1759
rect 151 -1766 159 -1759
rect 170 -1767 178 -1761
rect 255 -1777 265 -1767
rect 279 -1780 289 -1770
rect 368 -1767 375 -1761
rect 390 -1771 399 -1763
rect 434 -1770 442 -1763
rect 453 -1771 461 -1765
rect 538 -1781 548 -1771
rect 562 -1784 572 -1774
rect 630 -1775 636 -1769
rect 649 -1778 655 -1772
rect 670 -1778 676 -1772
rect 690 -1778 696 -1772
rect 721 -1775 727 -1769
rect 739 -1777 746 -1771
<< polysilicon >>
rect -110 1050 -109 1077
rect -167 1035 -146 1039
rect -167 1012 -166 1035
rect -147 1012 -146 1035
rect -181 959 -180 975
rect -246 938 -229 941
rect -230 917 -229 938
rect -1034 811 -552 819
rect -1034 810 -892 811
rect -1141 799 -1115 804
rect -1262 786 -1257 798
rect -1141 798 -1132 799
rect -1242 790 -1132 798
rect -1118 790 -1115 799
rect -1033 797 -1008 799
rect -1033 791 -1007 797
rect -1242 786 -1115 790
rect -1141 784 -1115 786
rect -1017 716 -1007 791
rect -963 754 -956 757
rect -899 754 -892 810
rect -760 754 -753 757
rect -696 754 -689 757
rect -573 754 -566 811
rect -509 754 -502 757
rect -392 754 -385 787
rect -328 754 -321 757
rect -963 716 -956 739
rect -1017 708 -956 716
rect -963 669 -956 708
rect -899 669 -892 739
rect -760 669 -753 739
rect -696 669 -689 739
rect -573 669 -566 739
rect -509 669 -502 739
rect -392 669 -385 739
rect -328 669 -321 739
rect -963 610 -956 654
rect -899 649 -892 654
rect -760 610 -753 654
rect -696 625 -689 654
rect -573 650 -566 654
rect -509 626 -502 654
rect -392 650 -385 654
rect -963 603 -753 610
rect -328 607 -321 654
rect -1006 464 -524 472
rect -1006 463 -864 464
rect -1143 452 -1026 453
rect -1143 443 -1142 452
rect -1128 444 -1036 452
rect -1005 450 -980 452
rect -1005 444 -979 450
rect -1128 443 -1026 444
rect -1143 442 -1026 443
rect -989 369 -979 444
rect -935 407 -928 410
rect -871 407 -864 463
rect -732 407 -725 410
rect -668 407 -661 410
rect -545 407 -538 464
rect -481 407 -474 410
rect -364 407 -357 440
rect -300 407 -293 410
rect -935 369 -928 392
rect -989 361 -928 369
rect -935 322 -928 361
rect -871 322 -864 392
rect -732 322 -725 392
rect -668 322 -661 392
rect -545 322 -538 392
rect -481 322 -474 392
rect -364 322 -357 392
rect -300 322 -293 392
rect -935 263 -928 307
rect -871 302 -864 307
rect -732 263 -725 307
rect -668 278 -661 307
rect -545 303 -538 307
rect -481 279 -474 307
rect -364 303 -357 307
rect -935 256 -725 263
rect -300 260 -293 307
rect -1006 78 -524 86
rect -1006 77 -864 78
rect -1190 64 -980 66
rect -1190 56 -979 64
rect -989 -17 -979 56
rect -935 21 -928 24
rect -871 21 -864 77
rect -732 21 -725 24
rect -668 21 -661 24
rect -545 21 -538 78
rect -481 21 -474 24
rect -364 21 -357 54
rect -300 21 -293 24
rect -935 -17 -928 6
rect -989 -25 -928 -17
rect -935 -64 -928 -25
rect -871 -64 -864 6
rect -732 -64 -725 6
rect -668 -64 -661 6
rect -545 -64 -538 6
rect -481 -64 -474 6
rect -364 -64 -357 6
rect -300 -64 -293 6
rect -935 -123 -928 -79
rect -871 -84 -864 -79
rect -732 -123 -725 -79
rect -668 -108 -661 -79
rect -545 -83 -538 -79
rect -481 -107 -474 -79
rect -364 -83 -357 -79
rect -935 -130 -725 -123
rect -300 -126 -293 -79
rect -1006 -346 -524 -338
rect -1006 -347 -864 -346
rect -1005 -360 -980 -358
rect -1005 -366 -979 -360
rect -989 -441 -979 -366
rect -935 -403 -928 -400
rect -871 -403 -864 -347
rect -732 -403 -725 -400
rect -668 -403 -661 -400
rect -545 -403 -538 -346
rect -481 -403 -474 -400
rect -364 -403 -357 -370
rect -300 -403 -293 -400
rect -935 -441 -928 -418
rect -989 -449 -928 -441
rect -935 -488 -928 -449
rect -871 -488 -864 -418
rect -732 -488 -725 -418
rect -668 -488 -661 -418
rect -545 -488 -538 -418
rect -481 -488 -474 -418
rect -364 -488 -357 -418
rect -300 -488 -293 -418
rect -935 -547 -928 -503
rect -871 -508 -864 -503
rect -732 -547 -725 -503
rect -668 -532 -661 -503
rect -545 -507 -538 -503
rect -481 -531 -474 -503
rect -364 -507 -357 -503
rect -935 -554 -725 -547
rect -300 -550 -293 -503
rect -246 -1431 -229 917
rect -200 -772 -180 959
rect -167 -230 -146 1012
rect -128 494 -109 1050
rect 195 539 542 540
rect 203 532 542 539
rect -128 481 17 494
rect 131 475 138 478
rect 195 475 202 528
rect 334 475 341 478
rect 398 475 405 478
rect 521 475 528 532
rect 935 526 950 534
rect 585 475 592 478
rect 702 475 709 508
rect 766 475 773 478
rect 871 469 878 472
rect 935 469 942 526
rect 1266 534 1722 536
rect 961 527 1722 534
rect 961 526 1282 527
rect 1074 469 1081 472
rect 1138 469 1145 472
rect 1261 469 1268 526
rect 1325 469 1332 472
rect 1442 469 1449 502
rect 1506 469 1513 472
rect 131 428 138 460
rect 131 390 138 417
rect 195 390 202 460
rect 334 390 341 460
rect 398 390 405 460
rect 521 394 528 460
rect 521 390 530 394
rect 585 390 592 460
rect 702 390 709 460
rect 766 390 773 460
rect 871 417 878 454
rect 871 384 878 408
rect 935 384 942 454
rect 1074 384 1081 454
rect 1138 384 1145 454
rect 1261 384 1268 454
rect 1325 384 1332 454
rect 1442 384 1449 454
rect 1506 384 1513 454
rect 131 331 138 375
rect 195 370 202 375
rect 334 331 341 375
rect 398 346 405 375
rect 131 324 341 331
rect 267 268 281 324
rect 521 284 530 375
rect 585 347 592 375
rect 702 371 709 375
rect 766 328 773 375
rect 871 325 878 369
rect 935 364 942 369
rect 1074 325 1081 369
rect 1138 340 1145 369
rect 1261 365 1268 369
rect 1325 341 1332 369
rect 1442 365 1449 369
rect 871 318 1081 325
rect 1506 322 1513 369
rect 432 274 538 284
rect 1655 277 1678 527
rect 268 261 280 268
rect -20 244 142 256
rect 278 250 280 261
rect 434 258 441 274
rect 521 267 530 274
rect 837 261 1680 277
rect 434 244 441 245
rect -20 136 -8 244
rect 838 224 847 261
rect 1655 255 1678 261
rect 95 215 847 224
rect 31 183 38 186
rect 95 183 103 215
rect 204 171 212 177
rect 314 179 321 182
rect 378 179 385 205
rect 31 136 38 168
rect -20 123 38 136
rect 31 98 38 123
rect 95 151 103 168
rect 95 98 102 151
rect 204 124 212 155
rect 170 123 212 124
rect 180 114 212 123
rect 204 93 212 114
rect 269 124 278 176
rect 487 167 495 173
rect 574 171 580 175
rect 615 171 621 175
rect 666 171 672 175
rect 314 125 321 164
rect 285 124 321 125
rect 269 116 321 124
rect 31 79 38 83
rect 95 78 102 83
rect 204 69 212 77
rect 231 48 239 114
rect 314 94 321 116
rect 378 94 385 164
rect 487 120 495 151
rect 453 119 495 120
rect 463 110 495 119
rect 574 110 580 160
rect 615 110 621 160
rect 666 138 672 160
rect 652 132 672 138
rect 666 110 672 132
rect 487 89 495 110
rect 314 75 321 79
rect 378 74 385 79
rect 487 65 495 73
rect 574 49 580 99
rect 527 48 581 49
rect 231 42 581 48
rect 232 41 581 42
rect 615 24 621 99
rect 666 94 672 99
rect 522 23 621 24
rect 534 15 621 23
rect 534 14 616 15
rect 252 -185 599 -184
rect 260 -192 599 -185
rect -172 -243 76 -230
rect -172 -245 93 -243
rect 188 -249 195 -246
rect 252 -249 259 -196
rect 391 -249 398 -246
rect 455 -249 462 -246
rect 578 -249 585 -192
rect 992 -198 1007 -190
rect 642 -249 649 -246
rect 759 -249 766 -216
rect 823 -249 830 -246
rect 928 -255 935 -252
rect 992 -255 999 -198
rect 1323 -190 1779 -188
rect 1018 -197 1779 -190
rect 1018 -198 1339 -197
rect 1131 -255 1138 -252
rect 1195 -255 1202 -252
rect 1318 -255 1325 -198
rect 1382 -255 1389 -252
rect 1499 -255 1506 -222
rect 1563 -255 1570 -252
rect 188 -296 195 -264
rect 188 -334 195 -307
rect 252 -334 259 -264
rect 391 -334 398 -264
rect 455 -334 462 -264
rect 578 -330 585 -264
rect 578 -334 587 -330
rect 642 -334 649 -264
rect 759 -334 766 -264
rect 823 -334 830 -264
rect 928 -307 935 -270
rect 928 -340 935 -316
rect 992 -340 999 -270
rect 1131 -340 1138 -270
rect 1195 -340 1202 -270
rect 1318 -340 1325 -270
rect 1382 -340 1389 -270
rect 1499 -340 1506 -270
rect 1563 -340 1570 -270
rect 188 -393 195 -349
rect 252 -354 259 -349
rect 391 -393 398 -349
rect 455 -378 462 -349
rect 188 -400 398 -393
rect 324 -456 338 -400
rect 578 -440 587 -349
rect 642 -377 649 -349
rect 759 -353 766 -349
rect 823 -396 830 -349
rect 928 -399 935 -355
rect 992 -360 999 -355
rect 1131 -399 1138 -355
rect 1195 -384 1202 -355
rect 1318 -359 1325 -355
rect 1382 -383 1389 -355
rect 1499 -359 1506 -355
rect 928 -406 1138 -399
rect 1563 -402 1570 -355
rect 489 -450 595 -440
rect 1712 -447 1735 -197
rect 325 -463 337 -456
rect 37 -480 199 -468
rect 335 -474 337 -463
rect 491 -466 498 -450
rect 578 -457 587 -450
rect 894 -463 1737 -447
rect 491 -480 498 -479
rect 37 -588 49 -480
rect 895 -500 904 -463
rect 1712 -469 1735 -463
rect 152 -509 904 -500
rect 88 -541 95 -538
rect 152 -541 160 -509
rect 261 -553 269 -547
rect 371 -545 378 -542
rect 435 -545 442 -519
rect 88 -588 95 -556
rect 37 -601 95 -588
rect 88 -626 95 -601
rect 152 -573 160 -556
rect 152 -626 159 -573
rect 261 -600 269 -569
rect 227 -601 269 -600
rect 237 -610 269 -601
rect 261 -631 269 -610
rect 326 -600 335 -548
rect 544 -557 552 -551
rect 631 -553 637 -549
rect 672 -553 678 -549
rect 723 -553 729 -549
rect 371 -599 378 -560
rect 342 -600 378 -599
rect 326 -608 378 -600
rect 88 -645 95 -641
rect 152 -646 159 -641
rect 261 -655 269 -647
rect 288 -676 296 -610
rect 371 -630 378 -608
rect 435 -630 442 -560
rect 544 -604 552 -573
rect 510 -605 552 -604
rect 520 -614 552 -605
rect 631 -614 637 -564
rect 672 -614 678 -564
rect 723 -586 729 -564
rect 709 -592 729 -586
rect 723 -614 729 -592
rect 544 -635 552 -614
rect 371 -649 378 -645
rect 435 -650 442 -645
rect 544 -659 552 -651
rect 631 -675 637 -625
rect 584 -676 638 -675
rect 288 -682 638 -676
rect 289 -683 638 -682
rect 672 -700 678 -625
rect 723 -630 729 -625
rect 579 -701 678 -700
rect 591 -709 678 -701
rect 591 -710 673 -709
rect -181 -791 -180 -772
rect 232 -775 579 -774
rect 240 -782 579 -775
rect -200 -794 -180 -791
rect 168 -839 175 -836
rect 232 -839 239 -786
rect 371 -839 378 -836
rect 435 -839 442 -836
rect 558 -839 565 -782
rect 972 -788 987 -780
rect 622 -839 629 -836
rect 739 -839 746 -806
rect 803 -839 810 -836
rect 908 -845 915 -842
rect 972 -845 979 -788
rect 1303 -780 1759 -778
rect 998 -787 1759 -780
rect 998 -788 1319 -787
rect 1111 -845 1118 -842
rect 1175 -845 1182 -842
rect 1298 -845 1305 -788
rect 1362 -845 1369 -842
rect 1479 -845 1486 -812
rect 1543 -845 1550 -842
rect 168 -886 175 -854
rect 168 -924 175 -897
rect 232 -924 239 -854
rect 371 -924 378 -854
rect 435 -924 442 -854
rect 558 -920 565 -854
rect 558 -924 567 -920
rect 622 -924 629 -854
rect 739 -924 746 -854
rect 803 -924 810 -854
rect 908 -897 915 -860
rect 908 -930 915 -906
rect 972 -930 979 -860
rect 1111 -930 1118 -860
rect 1175 -930 1182 -860
rect 1298 -930 1305 -860
rect 1362 -930 1369 -860
rect 1479 -930 1486 -860
rect 1543 -930 1550 -860
rect 168 -983 175 -939
rect 232 -944 239 -939
rect 371 -983 378 -939
rect 435 -968 442 -939
rect 168 -990 378 -983
rect 304 -1046 318 -990
rect 558 -1030 567 -939
rect 622 -967 629 -939
rect 739 -943 746 -939
rect 803 -986 810 -939
rect 908 -989 915 -945
rect 972 -950 979 -945
rect 1111 -989 1118 -945
rect 1175 -974 1182 -945
rect 1298 -949 1305 -945
rect 1362 -973 1369 -945
rect 1479 -949 1486 -945
rect 908 -996 1118 -989
rect 1543 -992 1550 -945
rect 469 -1040 575 -1030
rect 1692 -1037 1715 -787
rect 305 -1053 317 -1046
rect 17 -1070 179 -1058
rect 315 -1064 317 -1053
rect 471 -1056 478 -1040
rect 558 -1047 567 -1040
rect 874 -1053 1717 -1037
rect 471 -1070 478 -1069
rect 17 -1178 29 -1070
rect 875 -1090 884 -1053
rect 1692 -1059 1715 -1053
rect 132 -1099 884 -1090
rect 68 -1131 75 -1128
rect 132 -1131 140 -1099
rect 241 -1143 249 -1137
rect 351 -1135 358 -1132
rect 415 -1135 422 -1109
rect 68 -1178 75 -1146
rect 17 -1191 75 -1178
rect 68 -1216 75 -1191
rect 132 -1163 140 -1146
rect 132 -1216 139 -1163
rect 241 -1190 249 -1159
rect 207 -1191 249 -1190
rect 217 -1200 249 -1191
rect 241 -1221 249 -1200
rect 306 -1190 315 -1138
rect 524 -1147 532 -1141
rect 611 -1143 617 -1139
rect 652 -1143 658 -1139
rect 703 -1143 709 -1139
rect 351 -1189 358 -1150
rect 322 -1190 358 -1189
rect 306 -1198 358 -1190
rect 68 -1235 75 -1231
rect 132 -1236 139 -1231
rect 241 -1245 249 -1237
rect 268 -1266 276 -1200
rect 351 -1220 358 -1198
rect 415 -1220 422 -1150
rect 524 -1194 532 -1163
rect 490 -1195 532 -1194
rect 500 -1204 532 -1195
rect 611 -1204 617 -1154
rect 652 -1204 658 -1154
rect 703 -1176 709 -1154
rect 689 -1182 709 -1176
rect 703 -1204 709 -1182
rect 524 -1225 532 -1204
rect 351 -1239 358 -1235
rect 415 -1240 422 -1235
rect 524 -1249 532 -1241
rect 611 -1265 617 -1215
rect 564 -1266 618 -1265
rect 268 -1272 618 -1266
rect 269 -1273 618 -1272
rect 652 -1290 658 -1215
rect 703 -1220 709 -1215
rect 559 -1291 658 -1290
rect 571 -1299 658 -1291
rect 571 -1300 653 -1299
rect 260 -1399 607 -1398
rect 268 -1406 607 -1399
rect -244 -1444 -229 -1431
rect -244 -1457 -241 -1444
rect -230 -1457 -229 -1444
rect 196 -1463 203 -1460
rect 260 -1463 267 -1410
rect 399 -1463 406 -1460
rect 463 -1463 470 -1460
rect 586 -1463 593 -1406
rect 1000 -1412 1015 -1404
rect 650 -1463 657 -1460
rect 767 -1463 774 -1430
rect 831 -1463 838 -1460
rect 936 -1469 943 -1466
rect 1000 -1469 1007 -1412
rect 1331 -1404 1787 -1402
rect 1026 -1411 1787 -1404
rect 1026 -1412 1347 -1411
rect 1139 -1469 1146 -1466
rect 1203 -1469 1210 -1466
rect 1326 -1469 1333 -1412
rect 1390 -1469 1397 -1466
rect 1507 -1469 1514 -1436
rect 1571 -1469 1578 -1466
rect 196 -1510 203 -1478
rect 196 -1548 203 -1521
rect 260 -1548 267 -1478
rect 399 -1548 406 -1478
rect 463 -1548 470 -1478
rect 586 -1544 593 -1478
rect 586 -1548 595 -1544
rect 650 -1548 657 -1478
rect 767 -1548 774 -1478
rect 831 -1548 838 -1478
rect 936 -1521 943 -1484
rect 936 -1554 943 -1530
rect 1000 -1554 1007 -1484
rect 1139 -1554 1146 -1484
rect 1203 -1554 1210 -1484
rect 1326 -1554 1333 -1484
rect 1390 -1554 1397 -1484
rect 1507 -1554 1514 -1484
rect 1571 -1554 1578 -1484
rect 196 -1607 203 -1563
rect 260 -1568 267 -1563
rect 399 -1607 406 -1563
rect 463 -1592 470 -1563
rect 196 -1614 406 -1607
rect 332 -1670 346 -1614
rect 586 -1654 595 -1563
rect 650 -1591 657 -1563
rect 767 -1567 774 -1563
rect 831 -1610 838 -1563
rect 936 -1613 943 -1569
rect 1000 -1574 1007 -1569
rect 1139 -1613 1146 -1569
rect 1203 -1598 1210 -1569
rect 1326 -1573 1333 -1569
rect 1390 -1597 1397 -1569
rect 1507 -1573 1514 -1569
rect 936 -1620 1146 -1613
rect 1571 -1616 1578 -1569
rect 497 -1664 603 -1654
rect 1720 -1661 1743 -1411
rect 333 -1677 345 -1670
rect 45 -1694 207 -1682
rect 343 -1688 345 -1677
rect 499 -1680 506 -1664
rect 586 -1671 595 -1664
rect 902 -1677 1745 -1661
rect 499 -1694 506 -1693
rect 45 -1802 57 -1694
rect 903 -1714 912 -1677
rect 1720 -1683 1743 -1677
rect 160 -1723 912 -1714
rect 96 -1755 103 -1752
rect 160 -1755 168 -1723
rect 269 -1767 277 -1761
rect 379 -1759 386 -1756
rect 443 -1759 450 -1733
rect 96 -1802 103 -1770
rect 45 -1815 103 -1802
rect 96 -1840 103 -1815
rect 160 -1787 168 -1770
rect 160 -1840 167 -1787
rect 269 -1814 277 -1783
rect 235 -1815 277 -1814
rect 245 -1824 277 -1815
rect 269 -1845 277 -1824
rect 334 -1814 343 -1762
rect 552 -1771 560 -1765
rect 639 -1767 645 -1763
rect 680 -1767 686 -1763
rect 731 -1767 737 -1763
rect 379 -1813 386 -1774
rect 350 -1814 386 -1813
rect 334 -1822 386 -1814
rect 96 -1859 103 -1855
rect 160 -1860 167 -1855
rect 269 -1869 277 -1861
rect 296 -1890 304 -1824
rect 379 -1844 386 -1822
rect 443 -1844 450 -1774
rect 552 -1818 560 -1787
rect 518 -1819 560 -1818
rect 528 -1828 560 -1819
rect 639 -1828 645 -1778
rect 680 -1828 686 -1778
rect 731 -1800 737 -1778
rect 717 -1806 737 -1800
rect 731 -1828 737 -1806
rect 552 -1849 560 -1828
rect 379 -1863 386 -1859
rect 443 -1864 450 -1859
rect 552 -1873 560 -1865
rect 639 -1889 645 -1839
rect 592 -1890 646 -1889
rect 296 -1896 646 -1890
rect 297 -1897 646 -1896
rect 680 -1914 686 -1839
rect 731 -1844 737 -1839
rect 587 -1915 686 -1914
rect 599 -1923 686 -1915
rect 599 -1924 681 -1923
<< polycontact >>
rect -133 1050 -110 1083
rect -166 1012 -147 1035
rect -203 959 -181 978
rect -246 917 -230 938
rect -1045 809 -1034 820
rect -1257 785 -1242 799
rect -1132 790 -1118 799
rect -1046 791 -1033 799
rect -392 787 -385 794
rect -696 617 -689 625
rect -509 618 -502 626
rect -328 600 -321 607
rect -1017 462 -1006 473
rect -1142 443 -1128 452
rect -1036 444 -1025 452
rect -1018 444 -1005 452
rect -364 440 -357 447
rect -668 270 -661 278
rect -481 271 -474 279
rect -300 253 -293 260
rect -1017 76 -1006 87
rect -1206 55 -1190 67
rect -364 54 -357 61
rect -668 -116 -661 -108
rect -481 -115 -474 -107
rect -300 -133 -293 -126
rect -1017 -348 -1006 -337
rect -1018 -366 -1005 -358
rect -364 -370 -357 -363
rect -668 -540 -661 -532
rect -481 -539 -474 -531
rect -300 -557 -293 -550
rect 194 528 203 539
rect 17 480 36 496
rect 702 508 709 515
rect 950 525 961 535
rect 1442 502 1449 509
rect 131 417 138 428
rect 870 408 879 417
rect 398 338 405 346
rect 585 339 592 347
rect 766 321 773 328
rect 1138 332 1145 340
rect 1325 333 1332 341
rect 1506 315 1513 322
rect 142 244 152 259
rect 268 250 278 261
rect 434 245 441 258
rect 378 205 385 211
rect 268 176 278 187
rect 169 113 180 123
rect 231 114 239 126
rect 452 109 463 119
rect 647 132 652 138
rect 522 11 534 23
rect 251 -196 260 -185
rect 76 -243 94 -230
rect 759 -216 766 -209
rect 1007 -199 1018 -189
rect 1499 -222 1506 -215
rect 188 -307 195 -296
rect 927 -316 936 -307
rect 455 -386 462 -378
rect 642 -385 649 -377
rect 823 -403 830 -396
rect 1195 -392 1202 -384
rect 1382 -391 1389 -383
rect 1563 -409 1570 -402
rect 199 -480 209 -465
rect 325 -474 335 -463
rect 491 -479 498 -466
rect 435 -519 442 -513
rect 325 -548 335 -537
rect 226 -611 237 -601
rect 288 -610 296 -598
rect 509 -615 520 -605
rect 704 -592 709 -586
rect 579 -713 591 -701
rect -203 -791 -181 -772
rect 231 -786 240 -775
rect 739 -806 746 -799
rect 987 -789 998 -779
rect 1479 -812 1486 -805
rect 168 -897 175 -886
rect 907 -906 916 -897
rect 435 -976 442 -968
rect 622 -975 629 -967
rect 803 -993 810 -986
rect 1175 -982 1182 -974
rect 1362 -981 1369 -973
rect 1543 -999 1550 -992
rect 179 -1070 189 -1055
rect 305 -1064 315 -1053
rect 471 -1069 478 -1056
rect 415 -1109 422 -1103
rect 305 -1138 315 -1127
rect 206 -1201 217 -1191
rect 268 -1200 276 -1188
rect 489 -1205 500 -1195
rect 684 -1182 689 -1176
rect 559 -1303 571 -1291
rect 259 -1410 268 -1399
rect -241 -1460 -230 -1444
rect 767 -1430 774 -1423
rect 1015 -1413 1026 -1403
rect 1507 -1436 1514 -1429
rect 196 -1521 203 -1510
rect 935 -1530 944 -1521
rect 463 -1600 470 -1592
rect 650 -1599 657 -1591
rect 831 -1617 838 -1610
rect 1203 -1606 1210 -1598
rect 1390 -1605 1397 -1597
rect 1571 -1623 1578 -1616
rect 207 -1694 217 -1679
rect 333 -1688 343 -1677
rect 499 -1693 506 -1680
rect 443 -1733 450 -1727
rect 333 -1762 343 -1751
rect 234 -1825 245 -1815
rect 296 -1824 304 -1812
rect 517 -1829 528 -1819
rect 712 -1806 717 -1800
rect 587 -1927 599 -1915
<< metal1 >>
rect -382 1055 -133 1079
rect -110 1055 -76 1079
rect -381 1035 -148 1036
rect -381 1012 -166 1035
rect -381 1011 -148 1012
rect -376 959 -203 975
rect -181 959 -180 975
rect -380 918 -246 936
rect -230 918 -228 936
rect -1108 849 -78 867
rect -1104 824 -1090 849
rect -1171 809 -1045 824
rect -1262 799 -1243 803
rect -1262 785 -1257 799
rect -1242 785 -1240 788
rect -1262 768 -1240 785
rect -1258 728 -1240 768
rect -1171 754 -1157 809
rect -1129 799 -1049 801
rect -1118 791 -1046 799
rect -643 794 -384 796
rect -1118 790 -1049 791
rect -1129 788 -1049 790
rect -999 783 -658 793
rect -643 787 -392 794
rect -385 787 -384 794
rect -643 786 -384 787
rect -908 772 -900 783
rect -705 772 -697 783
rect -974 766 -900 772
rect -1076 754 -1063 757
rect -1171 740 -1063 754
rect -974 752 -967 766
rect -908 750 -900 766
rect -1503 711 -1240 728
rect -1258 710 -1240 711
rect -1076 482 -1063 740
rect -771 766 -697 772
rect -771 752 -764 766
rect -952 711 -943 742
rect -705 750 -697 766
rect -889 721 -881 742
rect -890 711 -881 721
rect -952 708 -881 711
rect -749 711 -740 742
rect -686 711 -678 742
rect -749 710 -678 711
rect -642 710 -633 786
rect -518 772 -510 781
rect -337 772 -329 781
rect -584 766 -510 772
rect -584 752 -577 766
rect -518 750 -510 766
rect -952 703 -855 708
rect -749 703 -633 710
rect -403 766 -329 772
rect -403 752 -396 766
rect -562 711 -553 742
rect -337 750 -329 766
rect -499 711 -491 742
rect -562 710 -491 711
rect -381 711 -372 742
rect -318 711 -310 742
rect -381 710 -310 711
rect -298 710 -190 712
rect -562 703 -445 710
rect -381 703 -190 710
rect -889 699 -855 703
rect -953 675 -904 683
rect -975 638 -967 660
rect -953 666 -943 675
rect -912 668 -904 675
rect -889 667 -881 699
rect -866 626 -855 699
rect -686 701 -633 703
rect -499 701 -445 703
rect -750 675 -701 683
rect -772 638 -764 660
rect -750 666 -740 675
rect -709 668 -701 675
rect -686 667 -678 701
rect -563 675 -514 683
rect -585 638 -577 660
rect -563 666 -553 675
rect -522 668 -514 675
rect -499 667 -491 701
rect -866 625 -509 626
rect -866 617 -696 625
rect -689 618 -509 625
rect -502 618 -468 626
rect -689 617 -468 618
rect -866 615 -468 617
rect -457 607 -445 701
rect -318 701 -190 703
rect -382 675 -333 683
rect -404 638 -396 660
rect -382 666 -372 675
rect -341 668 -333 675
rect -318 667 -310 701
rect -298 700 -190 701
rect -457 600 -328 607
rect -321 600 -288 607
rect -457 597 -288 600
rect -212 539 -195 700
rect -97 561 -78 849
rect -97 560 28 561
rect -97 546 965 560
rect -212 528 194 539
rect -212 526 203 528
rect 949 535 962 546
rect -212 525 23 526
rect 949 525 950 535
rect 961 525 962 535
rect 451 515 710 517
rect 174 504 436 514
rect 451 508 702 515
rect 709 508 710 515
rect 1191 509 1450 511
rect 451 507 710 508
rect -1080 473 -1063 482
rect 36 481 83 494
rect 186 493 194 504
rect 389 493 397 504
rect -1080 472 -1024 473
rect -1080 462 -1017 472
rect -1214 452 -1172 453
rect -1259 443 -1142 452
rect -1214 442 -1172 443
rect -1080 88 -1064 462
rect 71 459 83 481
rect 120 487 194 493
rect 120 473 127 487
rect 186 471 194 487
rect -1025 444 -1018 452
rect -615 447 -356 449
rect -971 436 -630 446
rect -615 440 -364 447
rect -357 440 -356 447
rect -615 439 -356 440
rect -880 425 -872 436
rect -677 425 -669 436
rect -946 419 -872 425
rect -946 405 -939 419
rect -880 403 -872 419
rect -743 419 -669 425
rect -743 405 -736 419
rect -924 364 -915 395
rect -677 403 -669 419
rect -861 374 -853 395
rect -862 364 -853 374
rect -924 361 -853 364
rect -721 364 -712 395
rect -658 364 -650 395
rect -721 363 -650 364
rect -614 363 -605 439
rect -490 425 -482 434
rect -309 425 -301 434
rect -556 419 -482 425
rect -556 405 -549 419
rect -490 403 -482 419
rect -924 356 -827 361
rect -721 356 -605 363
rect -375 419 -301 425
rect 74 431 83 459
rect 323 487 397 493
rect 323 473 330 487
rect 142 432 151 463
rect 389 471 397 487
rect 205 442 213 463
rect 204 432 213 442
rect 74 428 138 431
rect 74 419 131 428
rect -375 405 -368 419
rect -534 364 -525 395
rect -309 403 -301 419
rect 142 429 213 432
rect 345 432 354 463
rect 408 432 416 463
rect 345 431 416 432
rect 452 431 461 507
rect 576 493 584 502
rect 757 493 765 502
rect 835 498 1176 508
rect 1191 502 1442 509
rect 1449 502 1450 509
rect 1191 501 1450 502
rect 510 487 584 493
rect 510 473 517 487
rect 576 471 584 487
rect 142 424 239 429
rect 345 424 461 431
rect 691 487 765 493
rect 926 487 934 498
rect 1129 487 1137 498
rect 691 473 698 487
rect 532 432 541 463
rect 757 471 765 487
rect 595 432 603 463
rect 532 431 603 432
rect 860 481 934 487
rect 713 432 722 463
rect 776 432 784 463
rect 860 467 867 481
rect 926 465 934 481
rect 713 431 784 432
rect 1063 481 1137 487
rect 1063 467 1070 481
rect 532 424 649 431
rect 713 424 807 431
rect 205 420 239 424
rect -471 364 -463 395
rect -534 363 -463 364
rect -353 364 -344 395
rect -290 364 -282 395
rect 141 396 190 404
rect -353 363 -282 364
rect -274 363 -52 366
rect -534 356 -417 363
rect -353 356 -52 363
rect 119 359 127 381
rect 141 387 151 396
rect 182 389 190 396
rect 205 388 213 420
rect -861 352 -827 356
rect -925 328 -876 336
rect -947 291 -939 313
rect -925 319 -915 328
rect -884 321 -876 328
rect -861 320 -853 352
rect -838 279 -827 352
rect -658 354 -605 356
rect -471 354 -417 356
rect -722 328 -673 336
rect -744 291 -736 313
rect -722 319 -712 328
rect -681 321 -673 328
rect -658 320 -650 354
rect -535 328 -486 336
rect -557 291 -549 313
rect -535 319 -525 328
rect -494 321 -486 328
rect -471 320 -463 354
rect -838 278 -481 279
rect -838 270 -668 278
rect -661 271 -481 278
rect -474 271 -440 279
rect -661 270 -440 271
rect -838 268 -440 270
rect -429 260 -417 354
rect -290 355 -52 356
rect -290 354 -262 355
rect -354 328 -305 336
rect -376 291 -368 313
rect -354 319 -344 328
rect -313 321 -305 328
rect -290 320 -282 354
rect -429 253 -300 260
rect -293 253 -260 260
rect -429 250 -260 253
rect -1083 86 -1030 88
rect -1083 76 -1017 86
rect -1083 73 -1030 76
rect -1258 56 -1206 67
rect -1081 -337 -1062 73
rect -615 61 -356 63
rect -971 50 -630 60
rect -615 54 -364 61
rect -357 54 -356 61
rect -615 53 -356 54
rect -880 39 -872 50
rect -677 39 -669 50
rect -946 33 -872 39
rect -946 19 -939 33
rect -880 17 -872 33
rect -743 33 -669 39
rect -743 19 -736 33
rect -924 -22 -915 9
rect -677 17 -669 33
rect -861 -12 -853 9
rect -862 -22 -853 -12
rect -924 -25 -853 -22
rect -721 -22 -712 9
rect -658 -22 -650 9
rect -721 -23 -650 -22
rect -614 -23 -605 53
rect -490 39 -482 48
rect -309 39 -301 48
rect -556 33 -482 39
rect -556 19 -549 33
rect -490 17 -482 33
rect -924 -30 -827 -25
rect -721 -30 -605 -23
rect -375 33 -301 39
rect -375 19 -368 33
rect -534 -22 -525 9
rect -309 17 -301 33
rect -471 -22 -463 9
rect -534 -23 -463 -22
rect -353 -22 -344 9
rect -290 -22 -282 9
rect -353 -23 -282 -22
rect -223 -23 -210 -22
rect -534 -30 -417 -23
rect -353 -30 -206 -23
rect -861 -34 -827 -30
rect -925 -58 -876 -50
rect -947 -95 -939 -73
rect -925 -67 -915 -58
rect -884 -65 -876 -58
rect -861 -66 -853 -34
rect -838 -107 -827 -34
rect -658 -32 -605 -30
rect -471 -32 -417 -30
rect -722 -58 -673 -50
rect -744 -95 -736 -73
rect -722 -67 -712 -58
rect -681 -65 -673 -58
rect -658 -66 -650 -32
rect -535 -58 -486 -50
rect -557 -95 -549 -73
rect -535 -67 -525 -58
rect -494 -65 -486 -58
rect -471 -66 -463 -32
rect -838 -108 -481 -107
rect -838 -116 -668 -108
rect -661 -115 -481 -108
rect -474 -115 -440 -107
rect -661 -116 -440 -115
rect -838 -118 -440 -116
rect -429 -126 -417 -32
rect -290 -31 -206 -30
rect -290 -32 -262 -31
rect -354 -58 -305 -50
rect -376 -95 -368 -73
rect -354 -67 -344 -58
rect -313 -65 -305 -58
rect -290 -66 -282 -32
rect -429 -133 -300 -126
rect -293 -133 -260 -126
rect -429 -136 -260 -133
rect -1081 -338 -1028 -337
rect -1081 -348 -1017 -338
rect -1081 -349 -1028 -348
rect -1050 -351 -1028 -349
rect -1036 -366 -1018 -358
rect -615 -363 -356 -361
rect -971 -374 -630 -364
rect -615 -370 -364 -363
rect -357 -370 -356 -363
rect -615 -371 -356 -370
rect -880 -385 -872 -374
rect -677 -385 -669 -374
rect -946 -391 -872 -385
rect -946 -405 -939 -391
rect -880 -407 -872 -391
rect -743 -391 -669 -385
rect -743 -405 -736 -391
rect -924 -446 -915 -415
rect -677 -407 -669 -391
rect -861 -436 -853 -415
rect -862 -446 -853 -436
rect -924 -449 -853 -446
rect -721 -446 -712 -415
rect -658 -446 -650 -415
rect -721 -447 -650 -446
rect -614 -447 -605 -371
rect -490 -385 -482 -376
rect -309 -385 -301 -376
rect -556 -391 -482 -385
rect -556 -405 -549 -391
rect -490 -407 -482 -391
rect -924 -454 -827 -449
rect -721 -454 -605 -447
rect -375 -391 -301 -385
rect -375 -405 -368 -391
rect -534 -446 -525 -415
rect -309 -407 -301 -391
rect -471 -446 -463 -415
rect -534 -447 -463 -446
rect -353 -446 -344 -415
rect -290 -446 -282 -415
rect -353 -447 -282 -446
rect -271 -447 -258 -445
rect -534 -454 -417 -447
rect -353 -454 -258 -447
rect -861 -458 -827 -454
rect -925 -482 -876 -474
rect -947 -519 -939 -497
rect -925 -491 -915 -482
rect -884 -489 -876 -482
rect -861 -490 -853 -458
rect -838 -531 -827 -458
rect -658 -456 -605 -454
rect -471 -456 -417 -454
rect -722 -482 -673 -474
rect -744 -519 -736 -497
rect -722 -491 -712 -482
rect -681 -489 -673 -482
rect -658 -490 -650 -456
rect -535 -482 -486 -474
rect -557 -519 -549 -497
rect -535 -491 -525 -482
rect -494 -489 -486 -482
rect -471 -490 -463 -456
rect -838 -532 -481 -531
rect -838 -540 -668 -532
rect -661 -539 -481 -532
rect -474 -539 -440 -531
rect -661 -540 -440 -539
rect -838 -542 -440 -540
rect -429 -550 -417 -456
rect -290 -456 -258 -454
rect -354 -482 -305 -474
rect -376 -519 -368 -497
rect -354 -491 -344 -482
rect -313 -489 -305 -482
rect -290 -490 -282 -456
rect -429 -557 -300 -550
rect -293 -557 -285 -550
rect -429 -560 -285 -557
rect -271 -1397 -258 -456
rect -223 -823 -210 -31
rect -70 -184 -53 355
rect 228 347 239 420
rect 408 422 461 424
rect 595 422 649 424
rect 344 396 393 404
rect 322 359 330 381
rect 344 387 354 396
rect 385 389 393 396
rect 408 388 416 422
rect 531 396 580 404
rect 509 359 517 381
rect 531 387 541 396
rect 572 389 580 396
rect 595 388 603 422
rect 228 346 585 347
rect 228 338 398 346
rect 405 339 585 346
rect 592 339 626 347
rect 405 338 626 339
rect 228 336 626 338
rect 637 328 649 422
rect 776 422 807 424
rect 712 396 761 404
rect 690 359 698 381
rect 712 387 722 396
rect 753 389 761 396
rect 776 388 784 422
rect 799 416 807 422
rect 882 426 891 457
rect 1129 465 1137 481
rect 945 436 953 457
rect 944 426 953 436
rect 882 423 953 426
rect 1085 426 1094 457
rect 1148 426 1156 457
rect 1085 425 1156 426
rect 1192 425 1201 501
rect 1316 487 1324 496
rect 1497 487 1505 496
rect 1250 481 1324 487
rect 1250 467 1257 481
rect 1316 465 1324 481
rect 882 418 979 423
rect 1085 418 1201 425
rect 1431 481 1505 487
rect 1431 467 1438 481
rect 1272 426 1281 457
rect 1497 465 1505 481
rect 1335 426 1343 457
rect 1272 425 1343 426
rect 1453 426 1462 457
rect 1516 426 1524 457
rect 1453 425 1524 426
rect 1272 418 1389 425
rect 1453 418 1722 425
rect 799 408 870 416
rect 799 407 879 408
rect 945 414 979 418
rect 637 321 766 328
rect 773 321 806 328
rect 637 318 806 321
rect 821 300 834 407
rect 881 390 930 398
rect 859 353 867 375
rect 881 381 891 390
rect 922 383 930 390
rect 945 382 953 414
rect 968 341 979 414
rect 1148 416 1201 418
rect 1335 416 1389 418
rect 1084 390 1133 398
rect 1062 353 1070 375
rect 1084 381 1094 390
rect 1125 383 1133 390
rect 1148 382 1156 416
rect 1271 390 1320 398
rect 1249 353 1257 375
rect 1271 381 1281 390
rect 1312 383 1320 390
rect 1335 382 1343 416
rect 968 340 1325 341
rect 968 332 1138 340
rect 1145 333 1325 340
rect 1332 333 1366 341
rect 1145 332 1366 333
rect 968 330 1366 332
rect 1377 322 1389 416
rect 1516 417 1722 418
rect 1516 416 1535 417
rect 1702 416 1721 417
rect 1452 390 1501 398
rect 1430 353 1438 375
rect 1452 381 1462 390
rect 1493 383 1501 390
rect 1516 382 1524 416
rect 1564 382 1722 385
rect 1563 371 1722 382
rect 1563 369 1586 371
rect 1642 369 1722 371
rect 1377 315 1506 322
rect 1513 315 1546 322
rect 1377 312 1546 315
rect 140 288 837 300
rect 143 275 153 288
rect 1563 283 1579 369
rect 141 259 153 275
rect 1478 270 1619 283
rect 141 245 142 259
rect 152 245 153 259
rect 86 201 94 206
rect 20 195 94 201
rect 20 181 27 195
rect 86 179 94 195
rect 226 191 234 199
rect 191 185 234 191
rect 269 187 278 250
rect 434 211 441 245
rect 385 205 441 211
rect 369 197 377 202
rect 42 140 51 171
rect 191 171 199 185
rect 303 191 377 197
rect 303 177 310 191
rect 369 175 377 191
rect 509 187 517 195
rect 105 140 113 171
rect 42 138 113 140
rect 42 137 114 138
rect 42 132 139 137
rect 105 128 139 132
rect 41 104 90 112
rect 19 67 27 89
rect 41 95 51 104
rect 82 97 90 104
rect 105 96 113 128
rect 128 123 139 128
rect 214 125 224 158
rect 474 181 517 187
rect 325 136 334 167
rect 474 167 482 181
rect 565 179 588 185
rect 565 169 571 179
rect 388 136 396 167
rect 325 134 396 136
rect 656 169 662 185
rect 325 133 397 134
rect 325 128 422 133
rect 128 113 169 123
rect 214 116 231 125
rect 214 90 224 116
rect 239 116 241 125
rect 388 124 422 128
rect 324 100 373 108
rect 190 63 199 79
rect 302 63 310 85
rect 324 91 334 100
rect 365 93 373 100
rect 388 92 396 124
rect 411 119 422 124
rect 497 121 507 154
rect 584 147 590 160
rect 605 147 611 160
rect 584 141 611 147
rect 625 138 631 160
rect 674 140 681 161
rect 1478 140 1487 270
rect 625 132 647 138
rect 674 132 1487 140
rect 625 126 631 132
rect 411 109 452 119
rect 497 113 535 121
rect 584 120 631 126
rect 497 112 534 113
rect 497 86 507 112
rect 190 57 225 63
rect 473 59 482 75
rect 473 53 508 59
rect 523 23 534 112
rect 584 108 591 120
rect 624 108 631 120
rect 674 131 1478 132
rect 674 108 681 131
rect 565 88 571 102
rect 605 88 611 102
rect 565 83 634 88
rect 656 85 662 102
rect 751 -164 774 131
rect 76 -178 1022 -164
rect -72 -185 89 -184
rect -72 -196 251 -185
rect -72 -198 260 -196
rect 1006 -189 1019 -178
rect 12 -199 89 -198
rect 1006 -199 1007 -189
rect 1018 -199 1019 -189
rect 508 -209 767 -207
rect 231 -220 493 -210
rect 508 -216 759 -209
rect 766 -216 767 -209
rect 1248 -215 1507 -213
rect 508 -217 767 -216
rect 94 -243 140 -230
rect 243 -231 251 -220
rect 446 -231 454 -220
rect 128 -265 140 -243
rect 177 -237 251 -231
rect 177 -251 184 -237
rect 243 -253 251 -237
rect 131 -293 140 -265
rect 380 -237 454 -231
rect 380 -251 387 -237
rect 199 -292 208 -261
rect 446 -253 454 -237
rect 262 -282 270 -261
rect 261 -292 270 -282
rect 131 -296 195 -293
rect 131 -305 188 -296
rect 199 -295 270 -292
rect 402 -292 411 -261
rect 465 -292 473 -261
rect 402 -293 473 -292
rect 509 -293 518 -217
rect 633 -231 641 -222
rect 814 -231 822 -222
rect 892 -226 1233 -216
rect 1248 -222 1499 -215
rect 1506 -222 1507 -215
rect 1248 -223 1507 -222
rect 567 -237 641 -231
rect 567 -251 574 -237
rect 633 -253 641 -237
rect 199 -300 296 -295
rect 402 -300 518 -293
rect 748 -237 822 -231
rect 983 -237 991 -226
rect 1186 -237 1194 -226
rect 748 -251 755 -237
rect 589 -292 598 -261
rect 814 -253 822 -237
rect 652 -292 660 -261
rect 589 -293 660 -292
rect 917 -243 991 -237
rect 770 -292 779 -261
rect 833 -292 841 -261
rect 917 -257 924 -243
rect 983 -259 991 -243
rect 770 -293 841 -292
rect 1120 -243 1194 -237
rect 1120 -257 1127 -243
rect 589 -300 706 -293
rect 770 -300 864 -293
rect 262 -304 296 -300
rect 198 -328 247 -320
rect 176 -365 184 -343
rect 198 -337 208 -328
rect 239 -335 247 -328
rect 262 -336 270 -304
rect 285 -377 296 -304
rect 465 -302 518 -300
rect 652 -302 706 -300
rect 401 -328 450 -320
rect 379 -365 387 -343
rect 401 -337 411 -328
rect 442 -335 450 -328
rect 465 -336 473 -302
rect 588 -328 637 -320
rect 566 -365 574 -343
rect 588 -337 598 -328
rect 629 -335 637 -328
rect 652 -336 660 -302
rect 285 -378 642 -377
rect 285 -386 455 -378
rect 462 -385 642 -378
rect 649 -385 683 -377
rect 462 -386 683 -385
rect 285 -388 683 -386
rect 694 -396 706 -302
rect 833 -302 864 -300
rect 769 -328 818 -320
rect 747 -365 755 -343
rect 769 -337 779 -328
rect 810 -335 818 -328
rect 833 -336 841 -302
rect 856 -308 864 -302
rect 939 -298 948 -267
rect 1186 -259 1194 -243
rect 1002 -288 1010 -267
rect 1001 -298 1010 -288
rect 939 -301 1010 -298
rect 1142 -298 1151 -267
rect 1205 -298 1213 -267
rect 1142 -299 1213 -298
rect 1249 -299 1258 -223
rect 1373 -237 1381 -228
rect 1554 -237 1562 -228
rect 1307 -243 1381 -237
rect 1307 -257 1314 -243
rect 1373 -259 1381 -243
rect 939 -306 1036 -301
rect 1142 -306 1258 -299
rect 1488 -243 1562 -237
rect 1488 -257 1495 -243
rect 1329 -298 1338 -267
rect 1554 -259 1562 -243
rect 1392 -298 1400 -267
rect 1329 -299 1400 -298
rect 1510 -298 1519 -267
rect 1573 -298 1581 -267
rect 1510 -299 1581 -298
rect 1757 -299 1776 -298
rect 1329 -306 1446 -299
rect 1510 -306 1779 -299
rect 856 -316 927 -308
rect 856 -317 936 -316
rect 1002 -310 1036 -306
rect 694 -403 823 -396
rect 830 -403 863 -396
rect 694 -406 863 -403
rect 878 -424 891 -317
rect 938 -334 987 -326
rect 916 -371 924 -349
rect 938 -343 948 -334
rect 979 -341 987 -334
rect 1002 -342 1010 -310
rect 1025 -383 1036 -310
rect 1205 -308 1258 -306
rect 1392 -308 1446 -306
rect 1141 -334 1190 -326
rect 1119 -371 1127 -349
rect 1141 -343 1151 -334
rect 1182 -341 1190 -334
rect 1205 -342 1213 -308
rect 1328 -334 1377 -326
rect 1306 -371 1314 -349
rect 1328 -343 1338 -334
rect 1369 -341 1377 -334
rect 1392 -342 1400 -308
rect 1025 -384 1382 -383
rect 1025 -392 1195 -384
rect 1202 -391 1382 -384
rect 1389 -391 1423 -383
rect 1202 -392 1423 -391
rect 1025 -394 1423 -392
rect 1434 -402 1446 -308
rect 1573 -307 1779 -306
rect 1573 -308 1592 -307
rect 1509 -334 1558 -326
rect 1487 -371 1495 -349
rect 1509 -343 1519 -334
rect 1550 -341 1558 -334
rect 1573 -342 1581 -308
rect 1621 -342 1779 -339
rect 1620 -353 1779 -342
rect 1620 -355 1643 -353
rect 1699 -355 1779 -353
rect 1434 -409 1563 -402
rect 1570 -409 1603 -402
rect 1434 -412 1603 -409
rect 197 -436 894 -424
rect 200 -449 210 -436
rect 1620 -441 1636 -355
rect 198 -465 210 -449
rect 1535 -454 1676 -441
rect 198 -479 199 -465
rect 209 -479 210 -465
rect 143 -523 151 -518
rect 77 -529 151 -523
rect 77 -543 84 -529
rect 143 -545 151 -529
rect 283 -533 291 -525
rect 248 -539 291 -533
rect 326 -537 335 -474
rect 491 -513 498 -479
rect 442 -519 498 -513
rect 426 -527 434 -522
rect 99 -584 108 -553
rect 248 -553 256 -539
rect 360 -533 434 -527
rect 360 -547 367 -533
rect 426 -549 434 -533
rect 566 -537 574 -529
rect 162 -584 170 -553
rect 99 -586 170 -584
rect 99 -587 171 -586
rect 99 -592 196 -587
rect 162 -596 196 -592
rect 98 -620 147 -612
rect 76 -657 84 -635
rect 98 -629 108 -620
rect 139 -627 147 -620
rect 162 -628 170 -596
rect 185 -601 196 -596
rect 271 -599 281 -566
rect 531 -543 574 -537
rect 382 -588 391 -557
rect 531 -557 539 -543
rect 622 -545 645 -539
rect 622 -555 628 -545
rect 445 -588 453 -557
rect 382 -590 453 -588
rect 713 -555 719 -539
rect 382 -591 454 -590
rect 382 -596 479 -591
rect 185 -611 226 -601
rect 271 -608 288 -599
rect 271 -634 281 -608
rect 296 -608 298 -599
rect 445 -600 479 -596
rect 381 -624 430 -616
rect 247 -661 256 -645
rect 359 -661 367 -639
rect 381 -633 391 -624
rect 422 -631 430 -624
rect 445 -632 453 -600
rect 468 -605 479 -600
rect 554 -603 564 -570
rect 641 -577 647 -564
rect 662 -577 668 -564
rect 641 -583 668 -577
rect 682 -586 688 -564
rect 731 -584 738 -563
rect 1535 -584 1544 -454
rect 682 -592 704 -586
rect 731 -592 1544 -584
rect 682 -598 688 -592
rect 468 -615 509 -605
rect 554 -611 592 -603
rect 641 -604 688 -598
rect 554 -612 591 -611
rect 554 -638 564 -612
rect 247 -667 282 -661
rect 530 -665 539 -649
rect 530 -671 565 -665
rect 580 -701 591 -612
rect 641 -616 648 -604
rect 681 -616 688 -604
rect 731 -593 1535 -592
rect 731 -616 738 -593
rect 622 -636 628 -622
rect 662 -636 668 -622
rect 622 -641 691 -636
rect 713 -639 719 -622
rect 839 -754 852 -593
rect 56 -768 1002 -754
rect -181 -775 72 -774
rect -181 -786 231 -775
rect -181 -788 240 -786
rect 986 -779 999 -768
rect -181 -791 72 -788
rect 986 -789 987 -779
rect 998 -789 999 -779
rect 488 -799 747 -797
rect 211 -810 473 -800
rect 488 -806 739 -799
rect 746 -806 747 -799
rect 1228 -805 1487 -803
rect 488 -807 747 -806
rect 56 -823 120 -820
rect 223 -821 231 -810
rect 426 -821 434 -810
rect -223 -832 120 -823
rect -223 -833 66 -832
rect 73 -833 120 -832
rect -223 -842 -210 -833
rect 108 -855 120 -833
rect 157 -827 231 -821
rect 157 -841 164 -827
rect 223 -843 231 -827
rect 111 -883 120 -855
rect 360 -827 434 -821
rect 360 -841 367 -827
rect 179 -882 188 -851
rect 426 -843 434 -827
rect 242 -872 250 -851
rect 241 -882 250 -872
rect 111 -886 175 -883
rect 111 -895 168 -886
rect 179 -885 250 -882
rect 382 -882 391 -851
rect 445 -882 453 -851
rect 382 -883 453 -882
rect 489 -883 498 -807
rect 613 -821 621 -812
rect 794 -821 802 -812
rect 872 -816 1213 -806
rect 1228 -812 1479 -805
rect 1486 -812 1487 -805
rect 1228 -813 1487 -812
rect 547 -827 621 -821
rect 547 -841 554 -827
rect 613 -843 621 -827
rect 179 -890 276 -885
rect 382 -890 498 -883
rect 728 -827 802 -821
rect 963 -827 971 -816
rect 1166 -827 1174 -816
rect 728 -841 735 -827
rect 569 -882 578 -851
rect 794 -843 802 -827
rect 632 -882 640 -851
rect 569 -883 640 -882
rect 897 -833 971 -827
rect 750 -882 759 -851
rect 813 -882 821 -851
rect 897 -847 904 -833
rect 963 -849 971 -833
rect 750 -883 821 -882
rect 1100 -833 1174 -827
rect 1100 -847 1107 -833
rect 569 -890 686 -883
rect 750 -890 844 -883
rect 242 -894 276 -890
rect 178 -918 227 -910
rect 156 -955 164 -933
rect 178 -927 188 -918
rect 219 -925 227 -918
rect 242 -926 250 -894
rect 265 -967 276 -894
rect 445 -892 498 -890
rect 632 -892 686 -890
rect 381 -918 430 -910
rect 359 -955 367 -933
rect 381 -927 391 -918
rect 422 -925 430 -918
rect 445 -926 453 -892
rect 568 -918 617 -910
rect 546 -955 554 -933
rect 568 -927 578 -918
rect 609 -925 617 -918
rect 632 -926 640 -892
rect 265 -968 622 -967
rect 265 -976 435 -968
rect 442 -975 622 -968
rect 629 -975 663 -967
rect 442 -976 663 -975
rect 265 -978 663 -976
rect 674 -986 686 -892
rect 813 -892 844 -890
rect 749 -918 798 -910
rect 727 -955 735 -933
rect 749 -927 759 -918
rect 790 -925 798 -918
rect 813 -926 821 -892
rect 836 -898 844 -892
rect 919 -888 928 -857
rect 1166 -849 1174 -833
rect 982 -878 990 -857
rect 981 -888 990 -878
rect 919 -891 990 -888
rect 1122 -888 1131 -857
rect 1185 -888 1193 -857
rect 1122 -889 1193 -888
rect 1229 -889 1238 -813
rect 1353 -827 1361 -818
rect 1534 -827 1542 -818
rect 1287 -833 1361 -827
rect 1287 -847 1294 -833
rect 1353 -849 1361 -833
rect 919 -896 1016 -891
rect 1122 -896 1238 -889
rect 1468 -833 1542 -827
rect 1468 -847 1475 -833
rect 1309 -888 1318 -857
rect 1534 -849 1542 -833
rect 1372 -888 1380 -857
rect 1309 -889 1380 -888
rect 1490 -888 1499 -857
rect 1553 -888 1561 -857
rect 1490 -889 1561 -888
rect 1740 -889 1759 -888
rect 1309 -896 1426 -889
rect 1490 -896 1759 -889
rect 836 -906 907 -898
rect 836 -907 916 -906
rect 982 -900 1016 -896
rect 674 -993 803 -986
rect 810 -993 843 -986
rect 674 -996 843 -993
rect 858 -1014 871 -907
rect 918 -924 967 -916
rect 896 -961 904 -939
rect 918 -933 928 -924
rect 959 -931 967 -924
rect 982 -932 990 -900
rect 1005 -973 1016 -900
rect 1185 -898 1238 -896
rect 1372 -898 1426 -896
rect 1121 -924 1170 -916
rect 1099 -961 1107 -939
rect 1121 -933 1131 -924
rect 1162 -931 1170 -924
rect 1185 -932 1193 -898
rect 1308 -924 1357 -916
rect 1286 -961 1294 -939
rect 1308 -933 1318 -924
rect 1349 -931 1357 -924
rect 1372 -932 1380 -898
rect 1005 -974 1362 -973
rect 1005 -982 1175 -974
rect 1182 -981 1362 -974
rect 1369 -981 1403 -973
rect 1182 -982 1403 -981
rect 1005 -984 1403 -982
rect 1414 -992 1426 -898
rect 1553 -897 1759 -896
rect 1553 -898 1572 -897
rect 1489 -924 1538 -916
rect 1467 -961 1475 -939
rect 1489 -933 1499 -924
rect 1530 -931 1538 -924
rect 1553 -932 1561 -898
rect 1731 -929 1759 -928
rect 1601 -932 1759 -929
rect 1600 -943 1759 -932
rect 1600 -945 1623 -943
rect 1679 -945 1759 -943
rect 1414 -999 1543 -992
rect 1550 -999 1583 -992
rect 1414 -1002 1583 -999
rect 177 -1026 874 -1014
rect 180 -1039 190 -1026
rect 1600 -1031 1616 -945
rect 178 -1055 190 -1039
rect 1515 -1044 1656 -1031
rect 178 -1069 179 -1055
rect 189 -1069 190 -1055
rect 123 -1113 131 -1108
rect 57 -1119 131 -1113
rect 57 -1133 64 -1119
rect 123 -1135 131 -1119
rect 263 -1123 271 -1115
rect 228 -1129 271 -1123
rect 306 -1127 315 -1064
rect 471 -1103 478 -1069
rect 422 -1109 478 -1103
rect 406 -1117 414 -1112
rect 79 -1174 88 -1143
rect 228 -1143 236 -1129
rect 340 -1123 414 -1117
rect 340 -1137 347 -1123
rect 406 -1139 414 -1123
rect 546 -1127 554 -1119
rect 142 -1174 150 -1143
rect 79 -1176 150 -1174
rect 79 -1177 151 -1176
rect 79 -1182 176 -1177
rect 142 -1186 176 -1182
rect 78 -1210 127 -1202
rect 56 -1247 64 -1225
rect 78 -1219 88 -1210
rect 119 -1217 127 -1210
rect 142 -1218 150 -1186
rect 165 -1191 176 -1186
rect 251 -1189 261 -1156
rect 511 -1133 554 -1127
rect 362 -1178 371 -1147
rect 511 -1147 519 -1133
rect 602 -1135 625 -1129
rect 602 -1145 608 -1135
rect 425 -1178 433 -1147
rect 362 -1180 433 -1178
rect 693 -1145 699 -1129
rect 362 -1181 434 -1180
rect 362 -1186 459 -1181
rect 165 -1201 206 -1191
rect 251 -1198 268 -1189
rect 251 -1224 261 -1198
rect 276 -1198 278 -1189
rect 425 -1190 459 -1186
rect 361 -1214 410 -1206
rect 227 -1251 236 -1235
rect 339 -1251 347 -1229
rect 361 -1223 371 -1214
rect 402 -1221 410 -1214
rect 425 -1222 433 -1190
rect 448 -1195 459 -1190
rect 534 -1193 544 -1160
rect 621 -1167 627 -1154
rect 642 -1167 648 -1154
rect 621 -1173 648 -1167
rect 662 -1176 668 -1154
rect 711 -1174 718 -1153
rect 1515 -1174 1524 -1044
rect 662 -1182 684 -1176
rect 711 -1182 1524 -1174
rect 662 -1188 668 -1182
rect 448 -1205 489 -1195
rect 534 -1201 572 -1193
rect 621 -1194 668 -1188
rect 534 -1202 571 -1201
rect 534 -1228 544 -1202
rect 227 -1257 262 -1251
rect 510 -1255 519 -1239
rect 510 -1261 545 -1255
rect 560 -1291 571 -1202
rect 621 -1206 628 -1194
rect 661 -1206 668 -1194
rect 711 -1183 1515 -1182
rect 711 -1206 718 -1183
rect 602 -1226 608 -1212
rect 642 -1226 648 -1212
rect 602 -1231 671 -1226
rect 693 -1229 699 -1212
rect 879 -1378 893 -1183
rect 84 -1392 1030 -1378
rect -274 -1399 96 -1397
rect -274 -1410 259 -1399
rect -274 -1412 268 -1410
rect 1014 -1403 1027 -1392
rect -274 -1413 96 -1412
rect 1014 -1413 1015 -1403
rect 1026 -1413 1027 -1403
rect 516 -1423 775 -1421
rect 239 -1434 501 -1424
rect 516 -1430 767 -1423
rect 774 -1430 775 -1423
rect 1256 -1429 1515 -1427
rect 516 -1431 775 -1430
rect -254 -1444 87 -1443
rect -254 -1457 -241 -1444
rect -230 -1456 148 -1444
rect 251 -1445 259 -1434
rect 454 -1445 462 -1434
rect -230 -1457 87 -1456
rect 101 -1457 148 -1456
rect 136 -1479 148 -1457
rect 185 -1451 259 -1445
rect 185 -1465 192 -1451
rect 251 -1467 259 -1451
rect 139 -1507 148 -1479
rect 388 -1451 462 -1445
rect 388 -1465 395 -1451
rect 207 -1506 216 -1475
rect 454 -1467 462 -1451
rect 270 -1496 278 -1475
rect 269 -1506 278 -1496
rect 139 -1510 203 -1507
rect 139 -1519 196 -1510
rect 207 -1509 278 -1506
rect 410 -1506 419 -1475
rect 473 -1506 481 -1475
rect 410 -1507 481 -1506
rect 517 -1507 526 -1431
rect 641 -1445 649 -1436
rect 822 -1445 830 -1436
rect 900 -1440 1241 -1430
rect 1256 -1436 1507 -1429
rect 1514 -1436 1515 -1429
rect 1256 -1437 1515 -1436
rect 575 -1451 649 -1445
rect 575 -1465 582 -1451
rect 641 -1467 649 -1451
rect 207 -1514 304 -1509
rect 410 -1514 526 -1507
rect 756 -1451 830 -1445
rect 991 -1451 999 -1440
rect 1194 -1451 1202 -1440
rect 756 -1465 763 -1451
rect 597 -1506 606 -1475
rect 822 -1467 830 -1451
rect 660 -1506 668 -1475
rect 597 -1507 668 -1506
rect 925 -1457 999 -1451
rect 778 -1506 787 -1475
rect 841 -1506 849 -1475
rect 925 -1471 932 -1457
rect 991 -1473 999 -1457
rect 778 -1507 849 -1506
rect 1128 -1457 1202 -1451
rect 1128 -1471 1135 -1457
rect 597 -1514 714 -1507
rect 778 -1514 872 -1507
rect 270 -1518 304 -1514
rect 206 -1542 255 -1534
rect 184 -1579 192 -1557
rect 206 -1551 216 -1542
rect 247 -1549 255 -1542
rect 270 -1550 278 -1518
rect 293 -1591 304 -1518
rect 473 -1516 526 -1514
rect 660 -1516 714 -1514
rect 409 -1542 458 -1534
rect 387 -1579 395 -1557
rect 409 -1551 419 -1542
rect 450 -1549 458 -1542
rect 473 -1550 481 -1516
rect 596 -1542 645 -1534
rect 574 -1579 582 -1557
rect 596 -1551 606 -1542
rect 637 -1549 645 -1542
rect 660 -1550 668 -1516
rect 293 -1592 650 -1591
rect 293 -1600 463 -1592
rect 470 -1599 650 -1592
rect 657 -1599 691 -1591
rect 470 -1600 691 -1599
rect 293 -1602 691 -1600
rect 702 -1610 714 -1516
rect 841 -1516 872 -1514
rect 777 -1542 826 -1534
rect 755 -1579 763 -1557
rect 777 -1551 787 -1542
rect 818 -1549 826 -1542
rect 841 -1550 849 -1516
rect 864 -1522 872 -1516
rect 947 -1512 956 -1481
rect 1194 -1473 1202 -1457
rect 1010 -1502 1018 -1481
rect 1009 -1512 1018 -1502
rect 947 -1515 1018 -1512
rect 1150 -1512 1159 -1481
rect 1213 -1512 1221 -1481
rect 1150 -1513 1221 -1512
rect 1257 -1513 1266 -1437
rect 1381 -1451 1389 -1442
rect 1562 -1451 1570 -1442
rect 1315 -1457 1389 -1451
rect 1315 -1471 1322 -1457
rect 1381 -1473 1389 -1457
rect 947 -1520 1044 -1515
rect 1150 -1520 1266 -1513
rect 1496 -1457 1570 -1451
rect 1496 -1471 1503 -1457
rect 1337 -1512 1346 -1481
rect 1562 -1473 1570 -1457
rect 1400 -1512 1408 -1481
rect 1337 -1513 1408 -1512
rect 1518 -1512 1527 -1481
rect 1581 -1512 1589 -1481
rect 1518 -1513 1589 -1512
rect 1337 -1520 1454 -1513
rect 1518 -1520 1787 -1513
rect 864 -1530 935 -1522
rect 864 -1531 944 -1530
rect 1010 -1524 1044 -1520
rect 702 -1617 831 -1610
rect 838 -1617 871 -1610
rect 702 -1620 871 -1617
rect 886 -1638 899 -1531
rect 946 -1548 995 -1540
rect 924 -1585 932 -1563
rect 946 -1557 956 -1548
rect 987 -1555 995 -1548
rect 1010 -1556 1018 -1524
rect 1033 -1597 1044 -1524
rect 1213 -1522 1266 -1520
rect 1400 -1522 1454 -1520
rect 1149 -1548 1198 -1540
rect 1127 -1585 1135 -1563
rect 1149 -1557 1159 -1548
rect 1190 -1555 1198 -1548
rect 1213 -1556 1221 -1522
rect 1336 -1548 1385 -1540
rect 1314 -1585 1322 -1563
rect 1336 -1557 1346 -1548
rect 1377 -1555 1385 -1548
rect 1400 -1556 1408 -1522
rect 1033 -1598 1390 -1597
rect 1033 -1606 1203 -1598
rect 1210 -1605 1390 -1598
rect 1397 -1605 1431 -1597
rect 1210 -1606 1431 -1605
rect 1033 -1608 1431 -1606
rect 1442 -1616 1454 -1522
rect 1581 -1521 1787 -1520
rect 1581 -1522 1600 -1521
rect 1517 -1548 1566 -1540
rect 1495 -1585 1503 -1563
rect 1517 -1557 1527 -1548
rect 1558 -1555 1566 -1548
rect 1581 -1556 1589 -1522
rect 1629 -1556 1787 -1553
rect 1628 -1567 1787 -1556
rect 1628 -1569 1651 -1567
rect 1707 -1569 1787 -1567
rect 1442 -1623 1571 -1616
rect 1578 -1623 1611 -1616
rect 1442 -1626 1611 -1623
rect 205 -1650 902 -1638
rect 208 -1663 218 -1650
rect 1628 -1655 1644 -1569
rect 206 -1679 218 -1663
rect 1543 -1668 1684 -1655
rect 206 -1693 207 -1679
rect 217 -1693 218 -1679
rect 151 -1737 159 -1732
rect 85 -1743 159 -1737
rect 85 -1757 92 -1743
rect 151 -1759 159 -1743
rect 291 -1747 299 -1739
rect 256 -1753 299 -1747
rect 334 -1751 343 -1688
rect 499 -1727 506 -1693
rect 450 -1733 506 -1727
rect 434 -1741 442 -1736
rect 107 -1798 116 -1767
rect 256 -1767 264 -1753
rect 368 -1747 442 -1741
rect 368 -1761 375 -1747
rect 434 -1763 442 -1747
rect 574 -1751 582 -1743
rect 170 -1798 178 -1767
rect 107 -1800 178 -1798
rect 107 -1801 179 -1800
rect 107 -1806 204 -1801
rect 170 -1810 204 -1806
rect 106 -1834 155 -1826
rect 84 -1871 92 -1849
rect 106 -1843 116 -1834
rect 147 -1841 155 -1834
rect 170 -1842 178 -1810
rect 193 -1815 204 -1810
rect 279 -1813 289 -1780
rect 539 -1757 582 -1751
rect 390 -1802 399 -1771
rect 539 -1771 547 -1757
rect 630 -1759 653 -1753
rect 630 -1769 636 -1759
rect 453 -1802 461 -1771
rect 390 -1804 461 -1802
rect 721 -1769 727 -1753
rect 390 -1805 462 -1804
rect 390 -1810 487 -1805
rect 193 -1825 234 -1815
rect 279 -1822 296 -1813
rect 279 -1848 289 -1822
rect 304 -1822 306 -1813
rect 453 -1814 487 -1810
rect 389 -1838 438 -1830
rect 255 -1875 264 -1859
rect 367 -1875 375 -1853
rect 389 -1847 399 -1838
rect 430 -1845 438 -1838
rect 453 -1846 461 -1814
rect 476 -1819 487 -1814
rect 562 -1817 572 -1784
rect 649 -1791 655 -1778
rect 670 -1791 676 -1778
rect 649 -1797 676 -1791
rect 690 -1800 696 -1778
rect 739 -1798 746 -1777
rect 1543 -1798 1552 -1668
rect 690 -1806 712 -1800
rect 739 -1806 1552 -1798
rect 690 -1812 696 -1806
rect 476 -1829 517 -1819
rect 562 -1825 600 -1817
rect 649 -1818 696 -1812
rect 562 -1826 599 -1825
rect 562 -1852 572 -1826
rect 255 -1881 290 -1875
rect 538 -1879 547 -1863
rect 538 -1885 573 -1879
rect 588 -1915 599 -1826
rect 649 -1830 656 -1818
rect 689 -1830 696 -1818
rect 739 -1807 1543 -1806
rect 739 -1830 746 -1807
rect 630 -1850 636 -1836
rect 670 -1850 676 -1836
rect 630 -1855 699 -1850
rect 721 -1853 727 -1836
<< labels >>
rlabel metal1 125 363 126 367 1 gnd
rlabel metal1 158 488 159 492 5 vdd
rlabel metal1 328 363 329 367 1 gnd
rlabel metal1 361 488 362 492 5 vdd
rlabel metal1 515 363 516 367 1 gnd
rlabel metal1 548 488 549 492 5 vdd
rlabel metal1 696 363 697 367 1 gnd
rlabel metal1 729 488 730 492 5 vdd
rlabel metal1 865 357 866 361 1 gnd
rlabel metal1 898 482 899 486 5 vdd
rlabel metal1 1068 357 1069 361 1 gnd
rlabel metal1 1101 482 1102 486 5 vdd
rlabel metal1 1255 357 1256 361 1 gnd
rlabel metal1 1288 482 1289 486 5 vdd
rlabel metal1 1436 357 1437 361 1 gnd
rlabel metal1 1469 482 1470 486 5 vdd
rlabel metal1 209 188 211 190 5 vdd
rlabel metal1 219 59 221 61 1 gnd
rlabel metal1 58 196 59 200 5 vdd
rlabel metal1 25 71 26 75 1 gnd
rlabel metal1 492 184 494 186 5 vdd
rlabel metal1 502 55 504 57 1 gnd
rlabel metal1 341 192 342 196 5 vdd
rlabel metal1 308 67 309 71 1 gnd
rlabel metal1 569 182 570 183 5 vdd
rlabel metal1 568 86 569 87 1 gnd
rlabel metal1 658 90 659 92 1 gnd
rlabel metal1 658 180 659 182 5 vdd
rlabel metal1 -969 642 -968 646 1 gnd
rlabel metal1 -936 767 -935 771 5 vdd
rlabel metal1 -766 642 -765 646 1 gnd
rlabel metal1 -733 767 -732 771 5 vdd
rlabel metal1 -579 642 -578 646 1 gnd
rlabel metal1 -546 767 -545 771 5 vdd
rlabel metal1 -398 642 -397 646 1 gnd
rlabel metal1 -365 767 -364 771 5 vdd
rlabel metal1 -337 420 -336 424 5 vdd
rlabel metal1 -370 295 -369 299 1 gnd
rlabel metal1 -518 420 -517 424 5 vdd
rlabel metal1 -551 295 -550 299 1 gnd
rlabel metal1 -705 420 -704 424 5 vdd
rlabel metal1 -738 295 -737 299 1 gnd
rlabel metal1 -908 420 -907 424 5 vdd
rlabel metal1 -941 295 -940 299 1 gnd
rlabel metal1 -337 34 -336 38 5 vdd
rlabel metal1 -370 -91 -369 -87 1 gnd
rlabel metal1 -518 34 -517 38 5 vdd
rlabel metal1 -551 -91 -550 -87 1 gnd
rlabel metal1 -705 34 -704 38 5 vdd
rlabel metal1 -738 -91 -737 -87 1 gnd
rlabel metal1 -908 34 -907 38 5 vdd
rlabel metal1 -941 -91 -940 -87 1 gnd
rlabel metal1 -337 -390 -336 -386 5 vdd
rlabel metal1 -370 -515 -369 -511 1 gnd
rlabel metal1 -518 -390 -517 -386 5 vdd
rlabel metal1 -551 -515 -550 -511 1 gnd
rlabel metal1 -705 -390 -704 -386 5 vdd
rlabel metal1 -738 -515 -737 -511 1 gnd
rlabel metal1 -908 -390 -907 -386 5 vdd
rlabel metal1 -941 -515 -940 -511 1 gnd
rlabel metal1 182 -361 183 -357 1 gnd
rlabel metal1 215 -236 216 -232 5 vdd
rlabel metal1 385 -361 386 -357 1 gnd
rlabel metal1 418 -236 419 -232 5 vdd
rlabel metal1 572 -361 573 -357 1 gnd
rlabel metal1 605 -236 606 -232 5 vdd
rlabel metal1 753 -361 754 -357 1 gnd
rlabel metal1 786 -236 787 -232 5 vdd
rlabel metal1 922 -367 923 -363 1 gnd
rlabel metal1 955 -242 956 -238 5 vdd
rlabel metal1 1125 -367 1126 -363 1 gnd
rlabel metal1 1158 -242 1159 -238 5 vdd
rlabel metal1 1312 -367 1313 -363 1 gnd
rlabel metal1 1345 -242 1346 -238 5 vdd
rlabel metal1 1493 -367 1494 -363 1 gnd
rlabel metal1 1526 -242 1527 -238 5 vdd
rlabel metal1 266 -536 268 -534 5 vdd
rlabel metal1 276 -665 278 -663 1 gnd
rlabel metal1 115 -528 116 -524 5 vdd
rlabel metal1 82 -653 83 -649 1 gnd
rlabel metal1 549 -540 551 -538 5 vdd
rlabel metal1 559 -669 561 -667 1 gnd
rlabel metal1 398 -532 399 -528 5 vdd
rlabel metal1 365 -657 366 -653 1 gnd
rlabel metal1 626 -542 627 -541 5 vdd
rlabel metal1 625 -638 626 -637 1 gnd
rlabel metal1 715 -634 716 -632 1 gnd
rlabel metal1 715 -544 716 -542 5 vdd
rlabel metal1 162 -951 163 -947 1 gnd
rlabel metal1 195 -826 196 -822 5 vdd
rlabel metal1 365 -951 366 -947 1 gnd
rlabel metal1 398 -826 399 -822 5 vdd
rlabel metal1 552 -951 553 -947 1 gnd
rlabel metal1 585 -826 586 -822 5 vdd
rlabel metal1 733 -951 734 -947 1 gnd
rlabel metal1 766 -826 767 -822 5 vdd
rlabel metal1 902 -957 903 -953 1 gnd
rlabel metal1 935 -832 936 -828 5 vdd
rlabel metal1 1105 -957 1106 -953 1 gnd
rlabel metal1 1138 -832 1139 -828 5 vdd
rlabel metal1 1292 -957 1293 -953 1 gnd
rlabel metal1 1325 -832 1326 -828 5 vdd
rlabel metal1 1473 -957 1474 -953 1 gnd
rlabel metal1 1506 -832 1507 -828 5 vdd
rlabel metal1 246 -1126 248 -1124 5 vdd
rlabel metal1 256 -1255 258 -1253 1 gnd
rlabel metal1 95 -1118 96 -1114 5 vdd
rlabel metal1 62 -1243 63 -1239 1 gnd
rlabel metal1 529 -1130 531 -1128 5 vdd
rlabel metal1 539 -1259 541 -1257 1 gnd
rlabel metal1 378 -1122 379 -1118 5 vdd
rlabel metal1 345 -1247 346 -1243 1 gnd
rlabel metal1 606 -1132 607 -1131 5 vdd
rlabel metal1 605 -1228 606 -1227 1 gnd
rlabel metal1 695 -1224 696 -1222 1 gnd
rlabel metal1 695 -1134 696 -1132 5 vdd
rlabel metal1 190 -1575 191 -1571 1 gnd
rlabel metal1 223 -1450 224 -1446 5 vdd
rlabel metal1 393 -1575 394 -1571 1 gnd
rlabel metal1 426 -1450 427 -1446 5 vdd
rlabel metal1 580 -1575 581 -1571 1 gnd
rlabel metal1 613 -1450 614 -1446 5 vdd
rlabel metal1 761 -1575 762 -1571 1 gnd
rlabel metal1 794 -1450 795 -1446 5 vdd
rlabel metal1 930 -1581 931 -1577 1 gnd
rlabel metal1 963 -1456 964 -1452 5 vdd
rlabel metal1 1133 -1581 1134 -1577 1 gnd
rlabel metal1 1166 -1456 1167 -1452 5 vdd
rlabel metal1 1320 -1581 1321 -1577 1 gnd
rlabel metal1 1353 -1456 1354 -1452 5 vdd
rlabel metal1 1501 -1581 1502 -1577 1 gnd
rlabel metal1 1534 -1456 1535 -1452 5 vdd
rlabel metal1 274 -1750 276 -1748 5 vdd
rlabel metal1 284 -1879 286 -1877 1 gnd
rlabel metal1 123 -1742 124 -1738 5 vdd
rlabel metal1 90 -1867 91 -1863 1 gnd
rlabel metal1 557 -1754 559 -1752 5 vdd
rlabel metal1 567 -1883 569 -1881 1 gnd
rlabel metal1 406 -1746 407 -1742 5 vdd
rlabel metal1 373 -1871 374 -1867 1 gnd
rlabel metal1 634 -1756 635 -1755 5 vdd
rlabel metal1 633 -1852 634 -1851 1 gnd
rlabel metal1 723 -1848 724 -1846 1 gnd
rlabel metal1 723 -1758 724 -1756 5 vdd
<< end >>
