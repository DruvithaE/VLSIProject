magic
tech scmos
timestamp 1701500377
<< nwell >>
rect -674 5952 -543 5993
rect -471 5952 -340 5993
rect -284 5952 -153 5993
rect -103 5952 28 5993
rect 420 5673 551 5714
rect 623 5673 754 5714
rect 810 5673 941 5714
rect 991 5673 1122 5714
rect 1160 5667 1291 5708
rect 1363 5667 1494 5708
rect 1550 5667 1681 5708
rect 1731 5667 1862 5708
rect 2176 5665 2307 5706
rect 2345 5654 2411 5696
rect 3024 5687 3071 5712
rect -646 5605 -515 5646
rect -443 5605 -312 5646
rect -256 5605 -125 5646
rect -75 5605 56 5646
rect 3295 5610 3342 5635
rect 320 5381 451 5422
rect 489 5370 555 5412
rect 603 5377 734 5418
rect 772 5366 838 5408
rect 867 5381 955 5406
rect 961 5381 1014 5406
rect -646 5219 -515 5260
rect -443 5219 -312 5260
rect -256 5219 -125 5260
rect -75 5219 56 5260
rect 477 4949 608 4990
rect 680 4949 811 4990
rect 867 4949 998 4990
rect 1048 4949 1179 4990
rect 1217 4943 1348 4984
rect 1420 4943 1551 4984
rect 1607 4943 1738 4984
rect 1788 4943 1919 4984
rect 2174 4941 2305 4982
rect 2343 4930 2409 4972
rect -646 4795 -515 4836
rect -443 4795 -312 4836
rect -256 4795 -125 4836
rect -75 4795 56 4836
rect 377 4657 508 4698
rect 546 4646 612 4688
rect 660 4653 791 4694
rect 829 4642 895 4684
rect 924 4657 1012 4682
rect 1018 4657 1071 4682
rect 457 4359 588 4400
rect 660 4359 791 4400
rect 847 4359 978 4400
rect 1028 4359 1159 4400
rect 1197 4353 1328 4394
rect 1400 4353 1531 4394
rect 1587 4353 1718 4394
rect 1768 4353 1899 4394
rect 2175 4351 2306 4392
rect 2344 4340 2410 4382
rect 357 4067 488 4108
rect 526 4056 592 4098
rect 640 4063 771 4104
rect 809 4052 875 4094
rect 904 4067 992 4092
rect 998 4067 1051 4092
rect 485 3735 616 3776
rect 688 3735 819 3776
rect 875 3735 1006 3776
rect 1056 3735 1187 3776
rect 1225 3729 1356 3770
rect 1428 3729 1559 3770
rect 1615 3729 1746 3770
rect 1796 3729 1927 3770
rect 2176 3727 2307 3768
rect 2345 3716 2411 3758
rect 2178 3551 2309 3592
rect 2347 3540 2413 3582
rect 385 3443 516 3484
rect 554 3432 620 3474
rect 668 3439 799 3480
rect 837 3428 903 3470
rect 932 3443 1020 3468
rect 1026 3443 1079 3468
rect 527 2974 658 3015
rect 696 2963 762 3005
rect 444 2900 491 2925
rect 1494 2897 1714 2922
rect 527 2845 658 2846
rect 527 2805 721 2845
rect 751 2808 817 2850
rect 658 2804 721 2805
rect 2066 2765 2197 2806
rect 2203 2766 2265 2807
rect 2272 2772 2319 2797
rect 446 2738 493 2763
rect 507 2686 638 2687
rect 507 2685 696 2686
rect 507 2684 709 2685
rect 507 2646 764 2684
rect 771 2647 837 2689
rect 638 2645 764 2646
rect 702 2644 764 2645
rect 706 2643 764 2644
rect 445 2583 492 2608
rect 516 2467 647 2468
rect 516 2466 705 2467
rect 516 2465 718 2466
rect 516 2464 777 2465
rect 841 2464 907 2469
rect 516 2427 907 2464
rect 647 2426 843 2427
rect 711 2425 843 2426
rect 715 2424 843 2425
rect 774 2423 843 2424
rect 824 2422 843 2423
rect 445 2351 492 2376
rect 396 2037 527 2078
rect 599 2037 730 2078
rect 786 2037 917 2078
rect 967 2037 1098 2078
rect 1130 2033 1177 2058
rect 402 1748 533 1789
rect 605 1748 736 1789
rect 792 1748 923 1789
rect 973 1748 1104 1789
rect 1132 1741 1179 1766
rect 422 1431 553 1472
rect 625 1431 756 1472
rect 812 1431 943 1472
rect 993 1431 1124 1472
rect 1345 1463 1476 1504
rect 1482 1464 1613 1505
rect 1619 1460 1666 1485
rect 2066 1466 2197 1507
rect 2203 1467 2265 1508
rect 2272 1473 2319 1498
rect 1157 1424 1204 1449
rect 420 1140 551 1181
rect 623 1140 754 1181
rect 810 1140 941 1181
rect 991 1140 1122 1181
rect 1166 1133 1213 1158
rect 5034 1017 5213 1042
rect 4777 980 4956 1005
rect 4533 825 4712 850
rect 473 708 604 749
rect 642 697 708 739
rect 390 634 437 659
rect 1554 631 1774 656
rect 2066 635 2197 676
rect 2203 636 2265 677
rect 2272 642 2319 667
rect 5235 644 5323 669
rect 5329 644 5382 669
rect 473 579 604 580
rect 473 539 667 579
rect 697 542 763 584
rect 604 538 667 539
rect 392 472 439 497
rect 453 420 584 421
rect 453 419 642 420
rect 453 418 655 419
rect 453 380 710 418
rect 717 381 783 423
rect 584 379 710 380
rect 648 378 710 379
rect 652 377 710 378
rect 391 317 438 342
rect 462 201 593 202
rect 462 200 651 201
rect 462 199 664 200
rect 462 198 723 199
rect 787 198 853 203
rect 462 161 853 198
rect 593 160 789 161
rect 657 159 789 160
rect 661 158 789 159
rect 720 157 789 158
rect 770 156 789 157
rect 391 85 438 110
rect 679 -339 810 -298
rect 848 -350 914 -308
rect 1267 -382 1398 -341
rect 1404 -381 1466 -340
rect 1473 -375 1520 -350
rect 681 -537 812 -496
rect 850 -548 916 -506
rect 1267 -572 1398 -531
rect 1404 -571 1466 -530
rect 1473 -565 1520 -540
rect 681 -735 812 -694
rect 850 -746 916 -704
rect 1267 -778 1398 -737
rect 1404 -777 1466 -736
rect 1473 -771 1520 -746
rect 681 -930 812 -889
rect 850 -941 916 -899
rect 1267 -968 1398 -927
rect 1404 -967 1466 -926
rect 1473 -961 1520 -936
<< ntransistor >>
rect -648 5882 -641 5897
rect -584 5882 -577 5897
rect -445 5882 -438 5897
rect -381 5882 -374 5897
rect -258 5882 -251 5897
rect -194 5882 -187 5897
rect -77 5882 -70 5897
rect -13 5882 -6 5897
rect -620 5535 -613 5550
rect -556 5535 -549 5550
rect -417 5535 -410 5550
rect -353 5535 -346 5550
rect -230 5535 -223 5550
rect -166 5535 -159 5550
rect -49 5535 -42 5550
rect 15 5535 22 5550
rect -620 5149 -613 5164
rect -556 5149 -549 5164
rect -417 5149 -410 5164
rect -353 5149 -346 5164
rect -230 5149 -223 5164
rect -166 5149 -159 5164
rect -49 5149 -42 5164
rect 15 5149 22 5164
rect -620 4725 -613 4740
rect -556 4725 -549 4740
rect -417 4725 -410 4740
rect -353 4725 -346 4740
rect -230 4725 -223 4740
rect -166 4725 -159 4740
rect -49 4725 -42 4740
rect 15 4725 22 4740
rect 446 5603 453 5618
rect 510 5603 517 5618
rect 649 5603 656 5618
rect 713 5603 720 5618
rect 836 5603 845 5618
rect 900 5603 907 5618
rect 1017 5603 1024 5618
rect 1081 5603 1088 5618
rect 1186 5597 1193 5612
rect 1250 5597 1257 5612
rect 1389 5597 1396 5612
rect 1453 5597 1460 5612
rect 1576 5597 1583 5612
rect 1640 5597 1647 5612
rect 1757 5597 1764 5612
rect 1821 5597 1828 5612
rect 3042 5644 3048 5653
rect 2202 5595 2209 5610
rect 2266 5595 2273 5610
rect 2375 5589 2383 5605
rect 3313 5567 3319 5576
rect 346 5311 353 5326
rect 410 5311 417 5326
rect 519 5305 527 5321
rect 629 5307 636 5322
rect 693 5307 700 5322
rect 889 5327 895 5338
rect 930 5327 936 5338
rect 981 5327 987 5338
rect 802 5301 810 5317
rect 503 4879 510 4894
rect 567 4879 574 4894
rect 706 4879 713 4894
rect 770 4879 777 4894
rect 893 4879 902 4894
rect 957 4879 964 4894
rect 1074 4879 1081 4894
rect 1138 4879 1145 4894
rect 1243 4873 1250 4888
rect 1307 4873 1314 4888
rect 1446 4873 1453 4888
rect 1510 4873 1517 4888
rect 1633 4873 1640 4888
rect 1697 4873 1704 4888
rect 1814 4873 1821 4888
rect 1878 4873 1885 4888
rect 2200 4871 2207 4886
rect 2264 4871 2271 4886
rect 403 4587 410 4602
rect 467 4587 474 4602
rect 576 4581 584 4597
rect 686 4583 693 4598
rect 750 4583 757 4598
rect 946 4603 952 4614
rect 987 4603 993 4614
rect 1038 4603 1044 4614
rect 859 4577 867 4593
rect 2373 4865 2381 4881
rect 483 4289 490 4304
rect 547 4289 554 4304
rect 686 4289 693 4304
rect 750 4289 757 4304
rect 873 4289 882 4304
rect 937 4289 944 4304
rect 1054 4289 1061 4304
rect 1118 4289 1125 4304
rect 1223 4283 1230 4298
rect 1287 4283 1294 4298
rect 1426 4283 1433 4298
rect 1490 4283 1497 4298
rect 1613 4283 1620 4298
rect 1677 4283 1684 4298
rect 1794 4283 1801 4298
rect 1858 4283 1865 4298
rect 2201 4281 2208 4296
rect 2265 4281 2272 4296
rect 383 3997 390 4012
rect 447 3997 454 4012
rect 556 3991 564 4007
rect 666 3993 673 4008
rect 730 3993 737 4008
rect 926 4013 932 4024
rect 967 4013 973 4024
rect 1018 4013 1024 4024
rect 839 3987 847 4003
rect 2374 4275 2382 4291
rect 511 3665 518 3680
rect 575 3665 582 3680
rect 714 3665 721 3680
rect 778 3665 785 3680
rect 901 3665 910 3680
rect 965 3665 972 3680
rect 1082 3665 1089 3680
rect 1146 3665 1153 3680
rect 1251 3659 1258 3674
rect 1315 3659 1322 3674
rect 1454 3659 1461 3674
rect 1518 3659 1525 3674
rect 1641 3659 1648 3674
rect 1705 3659 1712 3674
rect 1822 3659 1829 3674
rect 1886 3659 1893 3674
rect 2202 3657 2209 3672
rect 2266 3657 2273 3672
rect 2375 3651 2383 3667
rect 2204 3481 2211 3496
rect 2268 3481 2275 3496
rect 411 3373 418 3388
rect 475 3373 482 3388
rect 584 3367 592 3383
rect 2377 3475 2385 3491
rect 694 3369 701 3384
rect 758 3369 765 3384
rect 954 3389 960 3400
rect 995 3389 1001 3400
rect 1046 3389 1052 3400
rect 867 3363 875 3379
rect 553 2904 560 2919
rect 617 2904 624 2919
rect 726 2898 734 2914
rect 462 2857 468 2866
rect 1516 2843 1522 2854
rect 1557 2843 1563 2854
rect 1596 2843 1602 2854
rect 1639 2843 1645 2854
rect 1681 2843 1687 2854
rect 553 2735 560 2750
rect 617 2735 624 2750
rect 680 2734 687 2749
rect 781 2743 789 2759
rect 464 2695 470 2704
rect 533 2576 540 2591
rect 597 2576 604 2591
rect 660 2575 667 2590
rect 728 2573 735 2588
rect 801 2582 809 2598
rect 463 2540 469 2549
rect 542 2357 549 2372
rect 606 2357 613 2372
rect 669 2356 676 2371
rect 737 2354 744 2369
rect 796 2353 803 2368
rect 871 2362 879 2378
rect 463 2308 469 2317
rect 1148 1990 1154 1999
rect 422 1967 429 1982
rect 486 1967 493 1982
rect 625 1967 632 1982
rect 689 1967 696 1982
rect 812 1967 819 1982
rect 876 1967 883 1982
rect 993 1967 1000 1982
rect 1057 1967 1064 1982
rect 1150 1698 1156 1707
rect 428 1678 435 1693
rect 492 1678 499 1693
rect 631 1678 638 1693
rect 695 1678 702 1693
rect 818 1678 825 1693
rect 882 1678 889 1693
rect 999 1678 1006 1693
rect 1063 1678 1070 1693
rect 1175 1381 1181 1390
rect 448 1361 455 1376
rect 512 1361 519 1376
rect 651 1361 658 1376
rect 715 1361 722 1376
rect 838 1361 845 1376
rect 902 1361 909 1376
rect 1019 1361 1026 1376
rect 1083 1361 1090 1376
rect 1184 1090 1190 1099
rect 446 1070 453 1085
rect 510 1070 517 1085
rect 649 1070 656 1085
rect 713 1070 720 1085
rect 836 1070 843 1085
rect 900 1070 907 1085
rect 1017 1070 1024 1085
rect 1081 1070 1088 1085
rect 499 638 506 653
rect 563 638 570 653
rect 672 632 680 648
rect 408 591 414 600
rect 499 469 506 484
rect 563 469 570 484
rect 626 468 633 483
rect 727 477 735 493
rect 2290 2729 2296 2738
rect 2092 2695 2099 2710
rect 2156 2695 2164 2710
rect 2229 2696 2237 2711
rect 1637 1417 1643 1426
rect 2290 1430 2296 1439
rect 1371 1393 1378 1408
rect 1435 1393 1442 1408
rect 1508 1394 1515 1409
rect 1572 1394 1579 1409
rect 2092 1396 2099 1411
rect 2156 1396 2163 1411
rect 2229 1397 2236 1412
rect 410 429 416 438
rect 479 310 486 325
rect 543 310 550 325
rect 606 309 613 324
rect 674 307 681 322
rect 747 316 755 332
rect 409 274 415 283
rect 488 91 495 106
rect 552 91 559 106
rect 615 90 622 105
rect 683 88 690 103
rect 742 87 749 102
rect 817 96 825 112
rect 5056 963 5062 974
rect 5097 963 5103 974
rect 5138 963 5144 974
rect 5180 963 5186 974
rect 4799 926 4805 937
rect 4840 926 4846 937
rect 4881 926 4887 937
rect 4923 926 4929 937
rect 4555 771 4561 782
rect 4596 771 4602 782
rect 4637 771 4643 782
rect 4679 771 4685 782
rect 1576 577 1582 588
rect 1617 577 1623 588
rect 1656 577 1662 588
rect 1699 577 1705 588
rect 1741 577 1747 588
rect 2290 599 2296 608
rect 409 42 415 51
rect 2092 565 2099 580
rect 2156 565 2163 580
rect 2229 566 2236 581
rect 705 -409 712 -394
rect 769 -409 776 -394
rect 878 -415 886 -399
rect 1491 -418 1497 -409
rect 1293 -452 1300 -437
rect 1357 -452 1364 -437
rect 1430 -451 1438 -436
rect 707 -607 714 -592
rect 771 -607 778 -592
rect 880 -613 888 -597
rect 1491 -608 1497 -599
rect 1293 -642 1300 -627
rect 1357 -642 1364 -627
rect 1430 -641 1437 -626
rect 707 -805 714 -790
rect 771 -805 778 -790
rect 880 -811 888 -795
rect 5257 590 5263 601
rect 5298 590 5304 601
rect 5349 590 5355 601
rect 1491 -814 1497 -805
rect 1293 -848 1300 -833
rect 1357 -848 1364 -833
rect 1430 -847 1438 -832
rect 707 -1000 714 -985
rect 771 -1000 778 -985
rect 880 -1006 888 -990
rect 1491 -1004 1497 -995
rect 1293 -1038 1300 -1023
rect 1357 -1038 1364 -1023
rect 1430 -1037 1437 -1022
<< ptransistor >>
rect -648 5967 -641 5982
rect -584 5967 -577 5982
rect -445 5967 -438 5982
rect -381 5967 -374 5982
rect -258 5967 -251 5982
rect -194 5967 -187 5982
rect -77 5967 -70 5982
rect -13 5967 -6 5982
rect -620 5620 -613 5635
rect -556 5620 -549 5635
rect -417 5620 -410 5635
rect -353 5620 -346 5635
rect -230 5620 -223 5635
rect -166 5620 -159 5635
rect -49 5620 -42 5635
rect 15 5620 22 5635
rect -620 5234 -613 5249
rect -556 5234 -549 5249
rect -417 5234 -410 5249
rect -353 5234 -346 5249
rect -230 5234 -223 5249
rect -166 5234 -159 5249
rect -49 5234 -42 5249
rect 15 5234 22 5249
rect -620 4810 -613 4825
rect -556 4810 -549 4825
rect -417 4810 -410 4825
rect -353 4810 -346 4825
rect -230 4810 -223 4825
rect -166 4810 -159 4825
rect -49 4810 -42 4825
rect 15 4810 22 4825
rect 446 5688 453 5703
rect 510 5688 517 5703
rect 649 5688 656 5703
rect 713 5688 720 5703
rect 836 5688 843 5703
rect 900 5688 907 5703
rect 1017 5688 1024 5703
rect 1081 5688 1088 5703
rect 1186 5682 1193 5697
rect 1250 5682 1257 5697
rect 1389 5682 1396 5697
rect 1453 5682 1460 5697
rect 1576 5682 1583 5697
rect 1640 5682 1647 5697
rect 1757 5682 1764 5697
rect 1821 5682 1828 5697
rect 2202 5680 2209 5695
rect 2266 5680 2273 5695
rect 2375 5667 2383 5683
rect 3042 5695 3048 5704
rect 3313 5618 3319 5627
rect 346 5396 353 5411
rect 410 5396 418 5411
rect 519 5383 527 5399
rect 629 5392 636 5407
rect 693 5392 700 5407
rect 802 5379 810 5395
rect 889 5388 895 5399
rect 930 5388 936 5399
rect 981 5388 987 5399
rect 503 4964 510 4979
rect 567 4964 574 4979
rect 706 4964 713 4979
rect 770 4964 777 4979
rect 893 4964 900 4979
rect 957 4964 964 4979
rect 1074 4964 1081 4979
rect 1138 4964 1145 4979
rect 1243 4958 1250 4973
rect 1307 4958 1314 4973
rect 1446 4958 1453 4973
rect 1510 4958 1517 4973
rect 1633 4958 1640 4973
rect 1697 4958 1704 4973
rect 1814 4958 1821 4973
rect 1878 4958 1885 4973
rect 2200 4956 2207 4971
rect 2264 4956 2271 4971
rect 2373 4943 2381 4959
rect 403 4672 410 4687
rect 467 4672 475 4687
rect 576 4659 584 4675
rect 686 4668 693 4683
rect 750 4668 757 4683
rect 859 4655 867 4671
rect 946 4664 952 4675
rect 987 4664 993 4675
rect 1038 4664 1044 4675
rect 483 4374 490 4389
rect 547 4374 554 4389
rect 686 4374 693 4389
rect 750 4374 757 4389
rect 873 4374 880 4389
rect 937 4374 944 4389
rect 1054 4374 1061 4389
rect 1118 4374 1125 4389
rect 1223 4368 1230 4383
rect 1287 4368 1294 4383
rect 1426 4368 1433 4383
rect 1490 4368 1497 4383
rect 1613 4368 1620 4383
rect 1677 4368 1684 4383
rect 1794 4368 1801 4383
rect 1858 4368 1865 4383
rect 2201 4366 2208 4381
rect 2265 4366 2272 4381
rect 2374 4353 2382 4369
rect 383 4082 390 4097
rect 447 4082 455 4097
rect 556 4069 564 4085
rect 666 4078 673 4093
rect 730 4078 737 4093
rect 839 4065 847 4081
rect 926 4074 932 4085
rect 967 4074 973 4085
rect 1018 4074 1024 4085
rect 511 3750 518 3765
rect 575 3750 582 3765
rect 714 3750 721 3765
rect 778 3750 785 3765
rect 901 3750 908 3765
rect 965 3750 972 3765
rect 1082 3750 1089 3765
rect 1146 3750 1153 3765
rect 1251 3744 1258 3759
rect 1315 3744 1322 3759
rect 1454 3744 1461 3759
rect 1518 3744 1525 3759
rect 1641 3744 1648 3759
rect 1705 3744 1712 3759
rect 1822 3744 1829 3759
rect 1886 3744 1893 3759
rect 2202 3742 2209 3757
rect 2266 3742 2273 3757
rect 2375 3729 2383 3745
rect 2204 3566 2211 3581
rect 2268 3566 2275 3581
rect 2377 3553 2385 3569
rect 411 3458 418 3473
rect 475 3458 483 3473
rect 584 3445 592 3461
rect 694 3454 701 3469
rect 758 3454 765 3469
rect 867 3441 875 3457
rect 954 3450 960 3461
rect 995 3450 1001 3461
rect 1046 3450 1052 3461
rect 553 2989 560 3004
rect 617 2989 624 3004
rect 726 2976 734 2992
rect 462 2908 468 2917
rect 1516 2904 1522 2915
rect 1557 2904 1563 2915
rect 1596 2904 1602 2915
rect 1639 2904 1645 2915
rect 1681 2904 1687 2915
rect 553 2820 560 2835
rect 617 2820 624 2835
rect 464 2746 470 2755
rect 680 2819 687 2834
rect 781 2821 789 2837
rect 533 2661 540 2676
rect 597 2661 604 2676
rect 463 2591 469 2600
rect 660 2660 667 2675
rect 728 2658 735 2673
rect 801 2660 809 2676
rect 542 2442 549 2457
rect 606 2442 613 2457
rect 669 2441 676 2456
rect 463 2359 469 2368
rect 737 2439 744 2454
rect 796 2438 803 2453
rect 871 2440 879 2456
rect 422 2052 429 2067
rect 486 2052 493 2067
rect 625 2052 632 2067
rect 689 2052 696 2067
rect 812 2052 819 2067
rect 876 2052 883 2067
rect 993 2052 1000 2067
rect 1057 2052 1064 2067
rect 1148 2041 1154 2050
rect 428 1763 435 1778
rect 492 1763 499 1778
rect 631 1763 638 1778
rect 695 1763 702 1778
rect 818 1763 825 1778
rect 882 1763 889 1778
rect 999 1763 1006 1778
rect 1063 1763 1070 1778
rect 1150 1749 1156 1758
rect 448 1446 455 1461
rect 512 1446 519 1461
rect 651 1446 658 1461
rect 715 1446 722 1461
rect 838 1446 845 1461
rect 902 1446 909 1461
rect 1019 1446 1026 1461
rect 1083 1446 1090 1461
rect 1175 1432 1181 1441
rect 446 1155 453 1170
rect 510 1155 517 1170
rect 649 1155 656 1170
rect 713 1155 720 1170
rect 836 1155 843 1170
rect 900 1155 907 1170
rect 1017 1155 1024 1170
rect 1081 1155 1088 1170
rect 1184 1141 1190 1150
rect 499 723 506 738
rect 563 723 570 738
rect 672 710 680 726
rect 408 642 414 651
rect 499 554 506 569
rect 563 554 570 569
rect 410 480 416 489
rect 626 553 633 568
rect 727 555 735 571
rect 2092 2780 2099 2795
rect 2156 2780 2164 2795
rect 2229 2781 2237 2796
rect 2290 2780 2296 2789
rect 1371 1478 1378 1493
rect 1435 1478 1442 1493
rect 1508 1479 1515 1494
rect 1572 1479 1579 1494
rect 2092 1481 2099 1496
rect 2156 1481 2163 1496
rect 2229 1482 2237 1497
rect 1637 1468 1643 1477
rect 2290 1481 2296 1490
rect 479 395 486 410
rect 543 395 550 410
rect 409 325 415 334
rect 606 394 613 409
rect 674 392 681 407
rect 747 394 755 410
rect 488 176 495 191
rect 552 176 559 191
rect 615 175 622 190
rect 409 93 415 102
rect 683 173 690 188
rect 742 172 749 187
rect 817 174 825 190
rect 5056 1024 5062 1035
rect 5097 1024 5103 1035
rect 5138 1024 5144 1035
rect 5180 1024 5186 1035
rect 4799 987 4805 998
rect 4840 987 4846 998
rect 4881 987 4887 998
rect 4923 987 4929 998
rect 4555 832 4561 843
rect 4596 832 4602 843
rect 4637 832 4643 843
rect 4679 832 4685 843
rect 2092 650 2099 665
rect 2156 650 2163 665
rect 2229 651 2237 666
rect 1576 638 1582 649
rect 1617 638 1623 649
rect 1656 638 1662 649
rect 1699 638 1705 649
rect 1741 638 1747 649
rect 2290 650 2296 659
rect 705 -324 712 -309
rect 769 -324 776 -309
rect 878 -337 886 -321
rect 1293 -367 1300 -352
rect 1357 -367 1364 -352
rect 1430 -366 1438 -351
rect 1491 -367 1497 -358
rect 707 -522 714 -507
rect 771 -522 778 -507
rect 880 -535 888 -519
rect 1293 -557 1300 -542
rect 1357 -557 1364 -542
rect 1430 -556 1438 -541
rect 1491 -557 1497 -548
rect 707 -720 714 -705
rect 771 -720 778 -705
rect 880 -733 888 -717
rect 1293 -763 1300 -748
rect 1357 -763 1364 -748
rect 1430 -762 1438 -747
rect 1491 -763 1497 -754
rect 5257 651 5263 662
rect 5298 651 5304 662
rect 5349 651 5355 662
rect 707 -915 714 -900
rect 771 -915 778 -900
rect 880 -928 888 -912
rect 1293 -953 1300 -938
rect 1357 -953 1364 -938
rect 1430 -952 1438 -937
rect 1491 -953 1497 -944
<< ndiffusion >>
rect -662 5895 -648 5897
rect -662 5888 -660 5895
rect -652 5888 -648 5895
rect -662 5882 -648 5888
rect -641 5894 -622 5897
rect -641 5885 -638 5894
rect -628 5885 -622 5894
rect -641 5882 -622 5885
rect -603 5896 -584 5897
rect -603 5888 -597 5896
rect -589 5888 -584 5896
rect -603 5882 -584 5888
rect -577 5895 -563 5897
rect -577 5887 -574 5895
rect -566 5887 -563 5895
rect -577 5882 -563 5887
rect -459 5895 -445 5897
rect -459 5888 -457 5895
rect -449 5888 -445 5895
rect -459 5882 -445 5888
rect -438 5894 -419 5897
rect -438 5885 -435 5894
rect -425 5885 -419 5894
rect -438 5882 -419 5885
rect -400 5896 -381 5897
rect -400 5888 -394 5896
rect -386 5888 -381 5896
rect -400 5882 -381 5888
rect -374 5895 -360 5897
rect -374 5887 -371 5895
rect -363 5887 -360 5895
rect -374 5882 -360 5887
rect -272 5895 -258 5897
rect -272 5888 -270 5895
rect -262 5888 -258 5895
rect -272 5882 -258 5888
rect -251 5894 -232 5897
rect -251 5885 -248 5894
rect -238 5885 -232 5894
rect -251 5882 -232 5885
rect -213 5896 -194 5897
rect -213 5888 -207 5896
rect -199 5888 -194 5896
rect -213 5882 -194 5888
rect -187 5895 -173 5897
rect -187 5887 -184 5895
rect -176 5887 -173 5895
rect -187 5882 -173 5887
rect -91 5895 -77 5897
rect -91 5888 -89 5895
rect -81 5888 -77 5895
rect -91 5882 -77 5888
rect -70 5894 -51 5897
rect -70 5885 -67 5894
rect -57 5885 -51 5894
rect -70 5882 -51 5885
rect -32 5896 -13 5897
rect -32 5888 -26 5896
rect -18 5888 -13 5896
rect -32 5882 -13 5888
rect -6 5895 8 5897
rect -6 5887 -3 5895
rect 5 5887 8 5895
rect -6 5882 8 5887
rect -634 5548 -620 5550
rect -634 5541 -632 5548
rect -624 5541 -620 5548
rect -634 5535 -620 5541
rect -613 5547 -594 5550
rect -613 5538 -610 5547
rect -600 5538 -594 5547
rect -613 5535 -594 5538
rect -575 5549 -556 5550
rect -575 5541 -569 5549
rect -561 5541 -556 5549
rect -575 5535 -556 5541
rect -549 5548 -535 5550
rect -549 5540 -546 5548
rect -538 5540 -535 5548
rect -549 5535 -535 5540
rect -431 5548 -417 5550
rect -431 5541 -429 5548
rect -421 5541 -417 5548
rect -431 5535 -417 5541
rect -410 5547 -391 5550
rect -410 5538 -407 5547
rect -397 5538 -391 5547
rect -410 5535 -391 5538
rect -372 5549 -353 5550
rect -372 5541 -366 5549
rect -358 5541 -353 5549
rect -372 5535 -353 5541
rect -346 5548 -332 5550
rect -346 5540 -343 5548
rect -335 5540 -332 5548
rect -346 5535 -332 5540
rect -244 5548 -230 5550
rect -244 5541 -242 5548
rect -234 5541 -230 5548
rect -244 5535 -230 5541
rect -223 5547 -204 5550
rect -223 5538 -220 5547
rect -210 5538 -204 5547
rect -223 5535 -204 5538
rect -185 5549 -166 5550
rect -185 5541 -179 5549
rect -171 5541 -166 5549
rect -185 5535 -166 5541
rect -159 5548 -145 5550
rect -159 5540 -156 5548
rect -148 5540 -145 5548
rect -159 5535 -145 5540
rect -63 5548 -49 5550
rect -63 5541 -61 5548
rect -53 5541 -49 5548
rect -63 5535 -49 5541
rect -42 5547 -23 5550
rect -42 5538 -39 5547
rect -29 5538 -23 5547
rect -42 5535 -23 5538
rect -4 5549 15 5550
rect -4 5541 2 5549
rect 10 5541 15 5549
rect -4 5535 15 5541
rect 22 5548 36 5550
rect 22 5540 25 5548
rect 33 5540 36 5548
rect 22 5535 36 5540
rect -634 5162 -620 5164
rect -634 5155 -632 5162
rect -624 5155 -620 5162
rect -634 5149 -620 5155
rect -613 5161 -594 5164
rect -613 5152 -610 5161
rect -600 5152 -594 5161
rect -613 5149 -594 5152
rect -575 5163 -556 5164
rect -575 5155 -569 5163
rect -561 5155 -556 5163
rect -575 5149 -556 5155
rect -549 5162 -535 5164
rect -549 5154 -546 5162
rect -538 5154 -535 5162
rect -549 5149 -535 5154
rect -431 5162 -417 5164
rect -431 5155 -429 5162
rect -421 5155 -417 5162
rect -431 5149 -417 5155
rect -410 5161 -391 5164
rect -410 5152 -407 5161
rect -397 5152 -391 5161
rect -410 5149 -391 5152
rect -372 5163 -353 5164
rect -372 5155 -366 5163
rect -358 5155 -353 5163
rect -372 5149 -353 5155
rect -346 5162 -332 5164
rect -346 5154 -343 5162
rect -335 5154 -332 5162
rect -346 5149 -332 5154
rect -244 5162 -230 5164
rect -244 5155 -242 5162
rect -234 5155 -230 5162
rect -244 5149 -230 5155
rect -223 5161 -204 5164
rect -223 5152 -220 5161
rect -210 5152 -204 5161
rect -223 5149 -204 5152
rect -185 5163 -166 5164
rect -185 5155 -179 5163
rect -171 5155 -166 5163
rect -185 5149 -166 5155
rect -159 5162 -145 5164
rect -159 5154 -156 5162
rect -148 5154 -145 5162
rect -159 5149 -145 5154
rect -63 5162 -49 5164
rect -63 5155 -61 5162
rect -53 5155 -49 5162
rect -63 5149 -49 5155
rect -42 5161 -23 5164
rect -42 5152 -39 5161
rect -29 5152 -23 5161
rect -42 5149 -23 5152
rect -4 5163 15 5164
rect -4 5155 2 5163
rect 10 5155 15 5163
rect -4 5149 15 5155
rect 22 5162 36 5164
rect 22 5154 25 5162
rect 33 5154 36 5162
rect 22 5149 36 5154
rect -634 4738 -620 4740
rect -634 4731 -632 4738
rect -624 4731 -620 4738
rect -634 4725 -620 4731
rect -613 4737 -594 4740
rect -613 4728 -610 4737
rect -600 4728 -594 4737
rect -613 4725 -594 4728
rect -575 4739 -556 4740
rect -575 4731 -569 4739
rect -561 4731 -556 4739
rect -575 4725 -556 4731
rect -549 4738 -535 4740
rect -549 4730 -546 4738
rect -538 4730 -535 4738
rect -549 4725 -535 4730
rect -431 4738 -417 4740
rect -431 4731 -429 4738
rect -421 4731 -417 4738
rect -431 4725 -417 4731
rect -410 4737 -391 4740
rect -410 4728 -407 4737
rect -397 4728 -391 4737
rect -410 4725 -391 4728
rect -372 4739 -353 4740
rect -372 4731 -366 4739
rect -358 4731 -353 4739
rect -372 4725 -353 4731
rect -346 4738 -332 4740
rect -346 4730 -343 4738
rect -335 4730 -332 4738
rect -346 4725 -332 4730
rect -244 4738 -230 4740
rect -244 4731 -242 4738
rect -234 4731 -230 4738
rect -244 4725 -230 4731
rect -223 4737 -204 4740
rect -223 4728 -220 4737
rect -210 4728 -204 4737
rect -223 4725 -204 4728
rect -185 4739 -166 4740
rect -185 4731 -179 4739
rect -171 4731 -166 4739
rect -185 4725 -166 4731
rect -159 4738 -145 4740
rect -159 4730 -156 4738
rect -148 4730 -145 4738
rect -159 4725 -145 4730
rect -63 4738 -49 4740
rect -63 4731 -61 4738
rect -53 4731 -49 4738
rect -63 4725 -49 4731
rect -42 4737 -23 4740
rect -42 4728 -39 4737
rect -29 4728 -23 4737
rect -42 4725 -23 4728
rect -4 4739 15 4740
rect -4 4731 2 4739
rect 10 4731 15 4739
rect -4 4725 15 4731
rect 22 4738 36 4740
rect 22 4730 25 4738
rect 33 4730 36 4738
rect 22 4725 36 4730
rect 432 5616 446 5618
rect 432 5609 434 5616
rect 442 5609 446 5616
rect 432 5603 446 5609
rect 453 5615 472 5618
rect 453 5606 456 5615
rect 466 5606 472 5615
rect 453 5603 472 5606
rect 491 5617 510 5618
rect 491 5609 497 5617
rect 505 5609 510 5617
rect 491 5603 510 5609
rect 517 5616 531 5618
rect 517 5608 520 5616
rect 528 5608 531 5616
rect 517 5603 531 5608
rect 635 5616 649 5618
rect 635 5609 637 5616
rect 645 5609 649 5616
rect 635 5603 649 5609
rect 656 5615 675 5618
rect 656 5606 659 5615
rect 669 5606 675 5615
rect 656 5603 675 5606
rect 694 5617 713 5618
rect 694 5609 700 5617
rect 708 5609 713 5617
rect 694 5603 713 5609
rect 720 5616 734 5618
rect 720 5608 723 5616
rect 731 5608 734 5616
rect 720 5603 734 5608
rect 822 5616 836 5618
rect 822 5609 824 5616
rect 832 5609 836 5616
rect 822 5603 836 5609
rect 845 5615 862 5618
rect 845 5606 846 5615
rect 856 5606 862 5615
rect 845 5603 862 5606
rect 881 5617 900 5618
rect 881 5609 887 5617
rect 895 5609 900 5617
rect 881 5603 900 5609
rect 907 5616 921 5618
rect 907 5608 910 5616
rect 918 5608 921 5616
rect 907 5603 921 5608
rect 1003 5616 1017 5618
rect 1003 5609 1005 5616
rect 1013 5609 1017 5616
rect 1003 5603 1017 5609
rect 1024 5615 1043 5618
rect 1024 5606 1027 5615
rect 1037 5606 1043 5615
rect 1024 5603 1043 5606
rect 1062 5617 1081 5618
rect 1062 5609 1068 5617
rect 1076 5609 1081 5617
rect 1062 5603 1081 5609
rect 1088 5616 1102 5618
rect 1088 5608 1091 5616
rect 1099 5608 1102 5616
rect 1088 5603 1102 5608
rect 1172 5610 1186 5612
rect 1172 5603 1174 5610
rect 1182 5603 1186 5610
rect 1172 5597 1186 5603
rect 1193 5609 1212 5612
rect 1193 5600 1196 5609
rect 1206 5600 1212 5609
rect 1193 5597 1212 5600
rect 1231 5611 1250 5612
rect 1231 5603 1237 5611
rect 1245 5603 1250 5611
rect 1231 5597 1250 5603
rect 1257 5610 1271 5612
rect 1257 5602 1260 5610
rect 1268 5602 1271 5610
rect 1257 5597 1271 5602
rect 1375 5610 1389 5612
rect 1375 5603 1377 5610
rect 1385 5603 1389 5610
rect 1375 5597 1389 5603
rect 1396 5609 1415 5612
rect 1396 5600 1399 5609
rect 1409 5600 1415 5609
rect 1396 5597 1415 5600
rect 1434 5611 1453 5612
rect 1434 5603 1440 5611
rect 1448 5603 1453 5611
rect 1434 5597 1453 5603
rect 1460 5610 1474 5612
rect 1460 5602 1463 5610
rect 1471 5602 1474 5610
rect 1460 5597 1474 5602
rect 1562 5610 1576 5612
rect 1562 5603 1564 5610
rect 1572 5603 1576 5610
rect 1562 5597 1576 5603
rect 1583 5609 1602 5612
rect 1583 5600 1586 5609
rect 1596 5600 1602 5609
rect 1583 5597 1602 5600
rect 1621 5611 1640 5612
rect 1621 5603 1627 5611
rect 1635 5603 1640 5611
rect 1621 5597 1640 5603
rect 1647 5610 1661 5612
rect 1647 5602 1650 5610
rect 1658 5602 1661 5610
rect 1647 5597 1661 5602
rect 1743 5610 1757 5612
rect 1743 5603 1745 5610
rect 1753 5603 1757 5610
rect 1743 5597 1757 5603
rect 1764 5609 1783 5612
rect 1764 5600 1767 5609
rect 1777 5600 1783 5609
rect 1764 5597 1783 5600
rect 1802 5611 1821 5612
rect 1802 5603 1808 5611
rect 1816 5603 1821 5611
rect 1802 5597 1821 5603
rect 1828 5610 1842 5612
rect 1828 5602 1831 5610
rect 1839 5602 1842 5610
rect 1828 5597 1842 5602
rect 3040 5644 3042 5653
rect 3048 5644 3050 5653
rect 3058 5644 3063 5653
rect 2188 5608 2202 5610
rect 2188 5601 2190 5608
rect 2198 5601 2202 5608
rect 2188 5595 2202 5601
rect 2209 5607 2228 5610
rect 2209 5598 2212 5607
rect 2222 5598 2228 5607
rect 2209 5595 2228 5598
rect 2247 5609 2266 5610
rect 2247 5601 2253 5609
rect 2261 5601 2266 5609
rect 2247 5595 2266 5601
rect 2273 5608 2287 5610
rect 2273 5600 2276 5608
rect 2284 5600 2287 5608
rect 2273 5595 2287 5600
rect 2358 5601 2375 5605
rect 2358 5591 2360 5601
rect 2370 5591 2375 5601
rect 2358 5589 2375 5591
rect 2383 5602 2398 5605
rect 2383 5592 2385 5602
rect 2395 5592 2398 5602
rect 2383 5589 2398 5592
rect 3311 5567 3313 5576
rect 3319 5567 3321 5576
rect 3329 5567 3334 5576
rect 332 5324 346 5326
rect 332 5317 334 5324
rect 342 5317 346 5324
rect 332 5311 346 5317
rect 353 5323 372 5326
rect 353 5314 356 5323
rect 366 5314 372 5323
rect 353 5311 372 5314
rect 391 5325 410 5326
rect 391 5317 397 5325
rect 405 5317 410 5325
rect 391 5311 410 5317
rect 417 5324 431 5326
rect 417 5316 420 5324
rect 428 5316 431 5324
rect 417 5311 431 5316
rect 502 5317 519 5321
rect 502 5307 504 5317
rect 514 5307 519 5317
rect 502 5305 519 5307
rect 527 5318 542 5321
rect 527 5308 529 5318
rect 539 5308 542 5318
rect 527 5305 542 5308
rect 615 5320 629 5322
rect 615 5313 617 5320
rect 625 5313 629 5320
rect 615 5307 629 5313
rect 636 5319 655 5322
rect 636 5310 639 5319
rect 649 5310 655 5319
rect 636 5307 655 5310
rect 674 5321 693 5322
rect 674 5313 680 5321
rect 688 5313 693 5321
rect 674 5307 693 5313
rect 700 5320 714 5322
rect 700 5312 703 5320
rect 711 5312 714 5320
rect 878 5335 889 5338
rect 878 5330 880 5335
rect 886 5330 889 5335
rect 878 5327 889 5330
rect 895 5336 911 5338
rect 895 5330 899 5336
rect 906 5330 911 5336
rect 895 5327 911 5330
rect 916 5335 930 5338
rect 916 5330 920 5335
rect 926 5330 930 5335
rect 916 5327 930 5330
rect 936 5336 949 5338
rect 936 5330 939 5336
rect 946 5330 949 5336
rect 936 5327 949 5330
rect 965 5335 981 5338
rect 965 5330 971 5335
rect 977 5330 981 5335
rect 965 5327 981 5330
rect 987 5336 998 5338
rect 987 5330 989 5336
rect 996 5330 998 5336
rect 987 5327 998 5330
rect 700 5307 714 5312
rect 785 5313 802 5317
rect 785 5303 787 5313
rect 797 5303 802 5313
rect 785 5301 802 5303
rect 810 5314 825 5317
rect 810 5304 812 5314
rect 822 5304 825 5314
rect 810 5301 825 5304
rect 489 4892 503 4894
rect 489 4885 491 4892
rect 499 4885 503 4892
rect 489 4879 503 4885
rect 510 4891 529 4894
rect 510 4882 513 4891
rect 523 4882 529 4891
rect 510 4879 529 4882
rect 548 4893 567 4894
rect 548 4885 554 4893
rect 562 4885 567 4893
rect 548 4879 567 4885
rect 574 4892 588 4894
rect 574 4884 577 4892
rect 585 4884 588 4892
rect 574 4879 588 4884
rect 692 4892 706 4894
rect 692 4885 694 4892
rect 702 4885 706 4892
rect 692 4879 706 4885
rect 713 4891 732 4894
rect 713 4882 716 4891
rect 726 4882 732 4891
rect 713 4879 732 4882
rect 751 4893 770 4894
rect 751 4885 757 4893
rect 765 4885 770 4893
rect 751 4879 770 4885
rect 777 4892 791 4894
rect 777 4884 780 4892
rect 788 4884 791 4892
rect 777 4879 791 4884
rect 879 4892 893 4894
rect 879 4885 881 4892
rect 889 4885 893 4892
rect 879 4879 893 4885
rect 902 4891 919 4894
rect 902 4882 903 4891
rect 913 4882 919 4891
rect 902 4879 919 4882
rect 938 4893 957 4894
rect 938 4885 944 4893
rect 952 4885 957 4893
rect 938 4879 957 4885
rect 964 4892 978 4894
rect 964 4884 967 4892
rect 975 4884 978 4892
rect 964 4879 978 4884
rect 1060 4892 1074 4894
rect 1060 4885 1062 4892
rect 1070 4885 1074 4892
rect 1060 4879 1074 4885
rect 1081 4891 1100 4894
rect 1081 4882 1084 4891
rect 1094 4882 1100 4891
rect 1081 4879 1100 4882
rect 1119 4893 1138 4894
rect 1119 4885 1125 4893
rect 1133 4885 1138 4893
rect 1119 4879 1138 4885
rect 1145 4892 1159 4894
rect 1145 4884 1148 4892
rect 1156 4884 1159 4892
rect 1145 4879 1159 4884
rect 1229 4886 1243 4888
rect 1229 4879 1231 4886
rect 1239 4879 1243 4886
rect 1229 4873 1243 4879
rect 1250 4885 1269 4888
rect 1250 4876 1253 4885
rect 1263 4876 1269 4885
rect 1250 4873 1269 4876
rect 1288 4887 1307 4888
rect 1288 4879 1294 4887
rect 1302 4879 1307 4887
rect 1288 4873 1307 4879
rect 1314 4886 1328 4888
rect 1314 4878 1317 4886
rect 1325 4878 1328 4886
rect 1314 4873 1328 4878
rect 1432 4886 1446 4888
rect 1432 4879 1434 4886
rect 1442 4879 1446 4886
rect 1432 4873 1446 4879
rect 1453 4885 1472 4888
rect 1453 4876 1456 4885
rect 1466 4876 1472 4885
rect 1453 4873 1472 4876
rect 1491 4887 1510 4888
rect 1491 4879 1497 4887
rect 1505 4879 1510 4887
rect 1491 4873 1510 4879
rect 1517 4886 1531 4888
rect 1517 4878 1520 4886
rect 1528 4878 1531 4886
rect 1517 4873 1531 4878
rect 1619 4886 1633 4888
rect 1619 4879 1621 4886
rect 1629 4879 1633 4886
rect 1619 4873 1633 4879
rect 1640 4885 1659 4888
rect 1640 4876 1643 4885
rect 1653 4876 1659 4885
rect 1640 4873 1659 4876
rect 1678 4887 1697 4888
rect 1678 4879 1684 4887
rect 1692 4879 1697 4887
rect 1678 4873 1697 4879
rect 1704 4886 1718 4888
rect 1704 4878 1707 4886
rect 1715 4878 1718 4886
rect 1704 4873 1718 4878
rect 1800 4886 1814 4888
rect 1800 4879 1802 4886
rect 1810 4879 1814 4886
rect 1800 4873 1814 4879
rect 1821 4885 1840 4888
rect 1821 4876 1824 4885
rect 1834 4876 1840 4885
rect 1821 4873 1840 4876
rect 1859 4887 1878 4888
rect 1859 4879 1865 4887
rect 1873 4879 1878 4887
rect 1859 4873 1878 4879
rect 1885 4886 1899 4888
rect 1885 4878 1888 4886
rect 1896 4878 1899 4886
rect 1885 4873 1899 4878
rect 2186 4884 2200 4886
rect 2186 4877 2188 4884
rect 2196 4877 2200 4884
rect 2186 4871 2200 4877
rect 2207 4883 2226 4886
rect 2207 4874 2210 4883
rect 2220 4874 2226 4883
rect 2207 4871 2226 4874
rect 2245 4885 2264 4886
rect 2245 4877 2251 4885
rect 2259 4877 2264 4885
rect 2245 4871 2264 4877
rect 2271 4884 2285 4886
rect 2271 4876 2274 4884
rect 2282 4876 2285 4884
rect 2271 4871 2285 4876
rect 2356 4877 2373 4881
rect 389 4600 403 4602
rect 389 4593 391 4600
rect 399 4593 403 4600
rect 389 4587 403 4593
rect 410 4599 429 4602
rect 410 4590 413 4599
rect 423 4590 429 4599
rect 410 4587 429 4590
rect 448 4601 467 4602
rect 448 4593 454 4601
rect 462 4593 467 4601
rect 448 4587 467 4593
rect 474 4600 488 4602
rect 474 4592 477 4600
rect 485 4592 488 4600
rect 474 4587 488 4592
rect 559 4593 576 4597
rect 559 4583 561 4593
rect 571 4583 576 4593
rect 559 4581 576 4583
rect 584 4594 599 4597
rect 584 4584 586 4594
rect 596 4584 599 4594
rect 584 4581 599 4584
rect 672 4596 686 4598
rect 672 4589 674 4596
rect 682 4589 686 4596
rect 672 4583 686 4589
rect 693 4595 712 4598
rect 693 4586 696 4595
rect 706 4586 712 4595
rect 693 4583 712 4586
rect 731 4597 750 4598
rect 731 4589 737 4597
rect 745 4589 750 4597
rect 731 4583 750 4589
rect 757 4596 771 4598
rect 757 4588 760 4596
rect 768 4588 771 4596
rect 935 4611 946 4614
rect 935 4606 937 4611
rect 943 4606 946 4611
rect 935 4603 946 4606
rect 952 4612 968 4614
rect 952 4606 956 4612
rect 963 4606 968 4612
rect 952 4603 968 4606
rect 973 4611 987 4614
rect 973 4606 977 4611
rect 983 4606 987 4611
rect 973 4603 987 4606
rect 993 4612 1006 4614
rect 993 4606 996 4612
rect 1003 4606 1006 4612
rect 993 4603 1006 4606
rect 1022 4611 1038 4614
rect 1022 4606 1028 4611
rect 1034 4606 1038 4611
rect 1022 4603 1038 4606
rect 1044 4612 1055 4614
rect 1044 4606 1046 4612
rect 1053 4606 1055 4612
rect 1044 4603 1055 4606
rect 757 4583 771 4588
rect 842 4589 859 4593
rect 842 4579 844 4589
rect 854 4579 859 4589
rect 842 4577 859 4579
rect 867 4590 882 4593
rect 867 4580 869 4590
rect 879 4580 882 4590
rect 867 4577 882 4580
rect 2356 4867 2358 4877
rect 2368 4867 2373 4877
rect 2356 4865 2373 4867
rect 2381 4878 2396 4881
rect 2381 4868 2383 4878
rect 2393 4868 2396 4878
rect 2381 4865 2396 4868
rect 469 4302 483 4304
rect 469 4295 471 4302
rect 479 4295 483 4302
rect 469 4289 483 4295
rect 490 4301 509 4304
rect 490 4292 493 4301
rect 503 4292 509 4301
rect 490 4289 509 4292
rect 528 4303 547 4304
rect 528 4295 534 4303
rect 542 4295 547 4303
rect 528 4289 547 4295
rect 554 4302 568 4304
rect 554 4294 557 4302
rect 565 4294 568 4302
rect 554 4289 568 4294
rect 672 4302 686 4304
rect 672 4295 674 4302
rect 682 4295 686 4302
rect 672 4289 686 4295
rect 693 4301 712 4304
rect 693 4292 696 4301
rect 706 4292 712 4301
rect 693 4289 712 4292
rect 731 4303 750 4304
rect 731 4295 737 4303
rect 745 4295 750 4303
rect 731 4289 750 4295
rect 757 4302 771 4304
rect 757 4294 760 4302
rect 768 4294 771 4302
rect 757 4289 771 4294
rect 859 4302 873 4304
rect 859 4295 861 4302
rect 869 4295 873 4302
rect 859 4289 873 4295
rect 882 4301 899 4304
rect 882 4292 883 4301
rect 893 4292 899 4301
rect 882 4289 899 4292
rect 918 4303 937 4304
rect 918 4295 924 4303
rect 932 4295 937 4303
rect 918 4289 937 4295
rect 944 4302 958 4304
rect 944 4294 947 4302
rect 955 4294 958 4302
rect 944 4289 958 4294
rect 1040 4302 1054 4304
rect 1040 4295 1042 4302
rect 1050 4295 1054 4302
rect 1040 4289 1054 4295
rect 1061 4301 1080 4304
rect 1061 4292 1064 4301
rect 1074 4292 1080 4301
rect 1061 4289 1080 4292
rect 1099 4303 1118 4304
rect 1099 4295 1105 4303
rect 1113 4295 1118 4303
rect 1099 4289 1118 4295
rect 1125 4302 1139 4304
rect 1125 4294 1128 4302
rect 1136 4294 1139 4302
rect 1125 4289 1139 4294
rect 1209 4296 1223 4298
rect 1209 4289 1211 4296
rect 1219 4289 1223 4296
rect 1209 4283 1223 4289
rect 1230 4295 1249 4298
rect 1230 4286 1233 4295
rect 1243 4286 1249 4295
rect 1230 4283 1249 4286
rect 1268 4297 1287 4298
rect 1268 4289 1274 4297
rect 1282 4289 1287 4297
rect 1268 4283 1287 4289
rect 1294 4296 1308 4298
rect 1294 4288 1297 4296
rect 1305 4288 1308 4296
rect 1294 4283 1308 4288
rect 1412 4296 1426 4298
rect 1412 4289 1414 4296
rect 1422 4289 1426 4296
rect 1412 4283 1426 4289
rect 1433 4295 1452 4298
rect 1433 4286 1436 4295
rect 1446 4286 1452 4295
rect 1433 4283 1452 4286
rect 1471 4297 1490 4298
rect 1471 4289 1477 4297
rect 1485 4289 1490 4297
rect 1471 4283 1490 4289
rect 1497 4296 1511 4298
rect 1497 4288 1500 4296
rect 1508 4288 1511 4296
rect 1497 4283 1511 4288
rect 1599 4296 1613 4298
rect 1599 4289 1601 4296
rect 1609 4289 1613 4296
rect 1599 4283 1613 4289
rect 1620 4295 1639 4298
rect 1620 4286 1623 4295
rect 1633 4286 1639 4295
rect 1620 4283 1639 4286
rect 1658 4297 1677 4298
rect 1658 4289 1664 4297
rect 1672 4289 1677 4297
rect 1658 4283 1677 4289
rect 1684 4296 1698 4298
rect 1684 4288 1687 4296
rect 1695 4288 1698 4296
rect 1684 4283 1698 4288
rect 1780 4296 1794 4298
rect 1780 4289 1782 4296
rect 1790 4289 1794 4296
rect 1780 4283 1794 4289
rect 1801 4295 1820 4298
rect 1801 4286 1804 4295
rect 1814 4286 1820 4295
rect 1801 4283 1820 4286
rect 1839 4297 1858 4298
rect 1839 4289 1845 4297
rect 1853 4289 1858 4297
rect 1839 4283 1858 4289
rect 1865 4296 1879 4298
rect 1865 4288 1868 4296
rect 1876 4288 1879 4296
rect 1865 4283 1879 4288
rect 2187 4294 2201 4296
rect 2187 4287 2189 4294
rect 2197 4287 2201 4294
rect 2187 4281 2201 4287
rect 2208 4293 2227 4296
rect 2208 4284 2211 4293
rect 2221 4284 2227 4293
rect 2208 4281 2227 4284
rect 2246 4295 2265 4296
rect 2246 4287 2252 4295
rect 2260 4287 2265 4295
rect 2246 4281 2265 4287
rect 2272 4294 2286 4296
rect 2272 4286 2275 4294
rect 2283 4286 2286 4294
rect 2272 4281 2286 4286
rect 2357 4287 2374 4291
rect 369 4010 383 4012
rect 369 4003 371 4010
rect 379 4003 383 4010
rect 369 3997 383 4003
rect 390 4009 409 4012
rect 390 4000 393 4009
rect 403 4000 409 4009
rect 390 3997 409 4000
rect 428 4011 447 4012
rect 428 4003 434 4011
rect 442 4003 447 4011
rect 428 3997 447 4003
rect 454 4010 468 4012
rect 454 4002 457 4010
rect 465 4002 468 4010
rect 454 3997 468 4002
rect 539 4003 556 4007
rect 539 3993 541 4003
rect 551 3993 556 4003
rect 539 3991 556 3993
rect 564 4004 579 4007
rect 564 3994 566 4004
rect 576 3994 579 4004
rect 564 3991 579 3994
rect 652 4006 666 4008
rect 652 3999 654 4006
rect 662 3999 666 4006
rect 652 3993 666 3999
rect 673 4005 692 4008
rect 673 3996 676 4005
rect 686 3996 692 4005
rect 673 3993 692 3996
rect 711 4007 730 4008
rect 711 3999 717 4007
rect 725 3999 730 4007
rect 711 3993 730 3999
rect 737 4006 751 4008
rect 737 3998 740 4006
rect 748 3998 751 4006
rect 915 4021 926 4024
rect 915 4016 917 4021
rect 923 4016 926 4021
rect 915 4013 926 4016
rect 932 4022 948 4024
rect 932 4016 936 4022
rect 943 4016 948 4022
rect 932 4013 948 4016
rect 953 4021 967 4024
rect 953 4016 957 4021
rect 963 4016 967 4021
rect 953 4013 967 4016
rect 973 4022 986 4024
rect 973 4016 976 4022
rect 983 4016 986 4022
rect 973 4013 986 4016
rect 1002 4021 1018 4024
rect 1002 4016 1008 4021
rect 1014 4016 1018 4021
rect 1002 4013 1018 4016
rect 1024 4022 1035 4024
rect 1024 4016 1026 4022
rect 1033 4016 1035 4022
rect 1024 4013 1035 4016
rect 737 3993 751 3998
rect 822 3999 839 4003
rect 822 3989 824 3999
rect 834 3989 839 3999
rect 822 3987 839 3989
rect 847 4000 862 4003
rect 847 3990 849 4000
rect 859 3990 862 4000
rect 847 3987 862 3990
rect 2357 4277 2359 4287
rect 2369 4277 2374 4287
rect 2357 4275 2374 4277
rect 2382 4288 2397 4291
rect 2382 4278 2384 4288
rect 2394 4278 2397 4288
rect 2382 4275 2397 4278
rect 497 3678 511 3680
rect 497 3671 499 3678
rect 507 3671 511 3678
rect 497 3665 511 3671
rect 518 3677 537 3680
rect 518 3668 521 3677
rect 531 3668 537 3677
rect 518 3665 537 3668
rect 556 3679 575 3680
rect 556 3671 562 3679
rect 570 3671 575 3679
rect 556 3665 575 3671
rect 582 3678 596 3680
rect 582 3670 585 3678
rect 593 3670 596 3678
rect 582 3665 596 3670
rect 700 3678 714 3680
rect 700 3671 702 3678
rect 710 3671 714 3678
rect 700 3665 714 3671
rect 721 3677 740 3680
rect 721 3668 724 3677
rect 734 3668 740 3677
rect 721 3665 740 3668
rect 759 3679 778 3680
rect 759 3671 765 3679
rect 773 3671 778 3679
rect 759 3665 778 3671
rect 785 3678 799 3680
rect 785 3670 788 3678
rect 796 3670 799 3678
rect 785 3665 799 3670
rect 887 3678 901 3680
rect 887 3671 889 3678
rect 897 3671 901 3678
rect 887 3665 901 3671
rect 910 3677 927 3680
rect 910 3668 911 3677
rect 921 3668 927 3677
rect 910 3665 927 3668
rect 946 3679 965 3680
rect 946 3671 952 3679
rect 960 3671 965 3679
rect 946 3665 965 3671
rect 972 3678 986 3680
rect 972 3670 975 3678
rect 983 3670 986 3678
rect 972 3665 986 3670
rect 1068 3678 1082 3680
rect 1068 3671 1070 3678
rect 1078 3671 1082 3678
rect 1068 3665 1082 3671
rect 1089 3677 1108 3680
rect 1089 3668 1092 3677
rect 1102 3668 1108 3677
rect 1089 3665 1108 3668
rect 1127 3679 1146 3680
rect 1127 3671 1133 3679
rect 1141 3671 1146 3679
rect 1127 3665 1146 3671
rect 1153 3678 1167 3680
rect 1153 3670 1156 3678
rect 1164 3670 1167 3678
rect 1153 3665 1167 3670
rect 1237 3672 1251 3674
rect 1237 3665 1239 3672
rect 1247 3665 1251 3672
rect 1237 3659 1251 3665
rect 1258 3671 1277 3674
rect 1258 3662 1261 3671
rect 1271 3662 1277 3671
rect 1258 3659 1277 3662
rect 1296 3673 1315 3674
rect 1296 3665 1302 3673
rect 1310 3665 1315 3673
rect 1296 3659 1315 3665
rect 1322 3672 1336 3674
rect 1322 3664 1325 3672
rect 1333 3664 1336 3672
rect 1322 3659 1336 3664
rect 1440 3672 1454 3674
rect 1440 3665 1442 3672
rect 1450 3665 1454 3672
rect 1440 3659 1454 3665
rect 1461 3671 1480 3674
rect 1461 3662 1464 3671
rect 1474 3662 1480 3671
rect 1461 3659 1480 3662
rect 1499 3673 1518 3674
rect 1499 3665 1505 3673
rect 1513 3665 1518 3673
rect 1499 3659 1518 3665
rect 1525 3672 1539 3674
rect 1525 3664 1528 3672
rect 1536 3664 1539 3672
rect 1525 3659 1539 3664
rect 1627 3672 1641 3674
rect 1627 3665 1629 3672
rect 1637 3665 1641 3672
rect 1627 3659 1641 3665
rect 1648 3671 1667 3674
rect 1648 3662 1651 3671
rect 1661 3662 1667 3671
rect 1648 3659 1667 3662
rect 1686 3673 1705 3674
rect 1686 3665 1692 3673
rect 1700 3665 1705 3673
rect 1686 3659 1705 3665
rect 1712 3672 1726 3674
rect 1712 3664 1715 3672
rect 1723 3664 1726 3672
rect 1712 3659 1726 3664
rect 1808 3672 1822 3674
rect 1808 3665 1810 3672
rect 1818 3665 1822 3672
rect 1808 3659 1822 3665
rect 1829 3671 1848 3674
rect 1829 3662 1832 3671
rect 1842 3662 1848 3671
rect 1829 3659 1848 3662
rect 1867 3673 1886 3674
rect 1867 3665 1873 3673
rect 1881 3665 1886 3673
rect 1867 3659 1886 3665
rect 1893 3672 1907 3674
rect 1893 3664 1896 3672
rect 1904 3664 1907 3672
rect 1893 3659 1907 3664
rect 2188 3670 2202 3672
rect 2188 3663 2190 3670
rect 2198 3663 2202 3670
rect 2188 3657 2202 3663
rect 2209 3669 2228 3672
rect 2209 3660 2212 3669
rect 2222 3660 2228 3669
rect 2209 3657 2228 3660
rect 2247 3671 2266 3672
rect 2247 3663 2253 3671
rect 2261 3663 2266 3671
rect 2247 3657 2266 3663
rect 2273 3670 2287 3672
rect 2273 3662 2276 3670
rect 2284 3662 2287 3670
rect 2273 3657 2287 3662
rect 2358 3663 2375 3667
rect 2358 3653 2360 3663
rect 2370 3653 2375 3663
rect 2358 3651 2375 3653
rect 2383 3664 2398 3667
rect 2383 3654 2385 3664
rect 2395 3654 2398 3664
rect 2383 3651 2398 3654
rect 2190 3494 2204 3496
rect 2190 3487 2192 3494
rect 2200 3487 2204 3494
rect 2190 3481 2204 3487
rect 2211 3493 2230 3496
rect 2211 3484 2214 3493
rect 2224 3484 2230 3493
rect 2211 3481 2230 3484
rect 2249 3495 2268 3496
rect 2249 3487 2255 3495
rect 2263 3487 2268 3495
rect 2249 3481 2268 3487
rect 2275 3494 2289 3496
rect 2275 3486 2278 3494
rect 2286 3486 2289 3494
rect 2275 3481 2289 3486
rect 2360 3487 2377 3491
rect 397 3386 411 3388
rect 397 3379 399 3386
rect 407 3379 411 3386
rect 397 3373 411 3379
rect 418 3385 437 3388
rect 418 3376 421 3385
rect 431 3376 437 3385
rect 418 3373 437 3376
rect 456 3387 475 3388
rect 456 3379 462 3387
rect 470 3379 475 3387
rect 456 3373 475 3379
rect 482 3386 496 3388
rect 482 3378 485 3386
rect 493 3378 496 3386
rect 482 3373 496 3378
rect 567 3379 584 3383
rect 567 3369 569 3379
rect 579 3369 584 3379
rect 567 3367 584 3369
rect 592 3380 607 3383
rect 592 3370 594 3380
rect 604 3370 607 3380
rect 592 3367 607 3370
rect 2360 3477 2362 3487
rect 2372 3477 2377 3487
rect 2360 3475 2377 3477
rect 2385 3488 2400 3491
rect 2385 3478 2387 3488
rect 2397 3478 2400 3488
rect 2385 3475 2400 3478
rect 680 3382 694 3384
rect 680 3375 682 3382
rect 690 3375 694 3382
rect 680 3369 694 3375
rect 701 3381 720 3384
rect 701 3372 704 3381
rect 714 3372 720 3381
rect 701 3369 720 3372
rect 739 3383 758 3384
rect 739 3375 745 3383
rect 753 3375 758 3383
rect 739 3369 758 3375
rect 765 3382 779 3384
rect 765 3374 768 3382
rect 776 3374 779 3382
rect 943 3397 954 3400
rect 943 3392 945 3397
rect 951 3392 954 3397
rect 943 3389 954 3392
rect 960 3398 976 3400
rect 960 3392 964 3398
rect 971 3392 976 3398
rect 960 3389 976 3392
rect 981 3397 995 3400
rect 981 3392 985 3397
rect 991 3392 995 3397
rect 981 3389 995 3392
rect 1001 3398 1014 3400
rect 1001 3392 1004 3398
rect 1011 3392 1014 3398
rect 1001 3389 1014 3392
rect 1030 3397 1046 3400
rect 1030 3392 1036 3397
rect 1042 3392 1046 3397
rect 1030 3389 1046 3392
rect 1052 3398 1063 3400
rect 1052 3392 1054 3398
rect 1061 3392 1063 3398
rect 1052 3389 1063 3392
rect 765 3369 779 3374
rect 850 3375 867 3379
rect 850 3365 852 3375
rect 862 3365 867 3375
rect 850 3363 867 3365
rect 875 3376 890 3379
rect 875 3366 877 3376
rect 887 3366 890 3376
rect 875 3363 890 3366
rect 539 2917 553 2919
rect 539 2910 541 2917
rect 549 2910 553 2917
rect 539 2904 553 2910
rect 560 2916 579 2919
rect 560 2907 563 2916
rect 573 2907 579 2916
rect 560 2904 579 2907
rect 598 2918 617 2919
rect 598 2910 604 2918
rect 612 2910 617 2918
rect 598 2904 617 2910
rect 624 2917 638 2919
rect 624 2909 627 2917
rect 635 2909 638 2917
rect 624 2904 638 2909
rect 709 2910 726 2914
rect 709 2900 711 2910
rect 721 2900 726 2910
rect 709 2898 726 2900
rect 734 2911 749 2914
rect 734 2901 736 2911
rect 746 2901 749 2911
rect 734 2898 749 2901
rect 460 2857 462 2866
rect 468 2857 470 2866
rect 478 2857 483 2866
rect 1505 2851 1516 2854
rect 1505 2846 1507 2851
rect 1513 2846 1516 2851
rect 1505 2843 1516 2846
rect 1522 2852 1538 2854
rect 1522 2846 1526 2852
rect 1533 2846 1538 2852
rect 1522 2843 1538 2846
rect 1543 2851 1557 2854
rect 1543 2846 1547 2851
rect 1553 2846 1557 2851
rect 1543 2843 1557 2846
rect 1563 2852 1576 2854
rect 1563 2846 1566 2852
rect 1573 2846 1576 2852
rect 1563 2843 1576 2846
rect 1582 2851 1596 2854
rect 1582 2845 1586 2851
rect 1592 2845 1596 2851
rect 1582 2843 1596 2845
rect 1602 2853 1615 2854
rect 1602 2846 1605 2853
rect 1612 2846 1615 2853
rect 1602 2843 1615 2846
rect 1625 2851 1639 2854
rect 1625 2845 1629 2851
rect 1635 2845 1639 2851
rect 1625 2843 1639 2845
rect 1645 2852 1658 2854
rect 1645 2846 1647 2852
rect 1654 2846 1658 2852
rect 1645 2843 1658 2846
rect 1665 2851 1681 2854
rect 1665 2846 1671 2851
rect 1677 2846 1681 2851
rect 1665 2843 1681 2846
rect 1687 2852 1698 2854
rect 1687 2846 1689 2852
rect 1696 2846 1698 2852
rect 1687 2843 1698 2846
rect 539 2748 553 2750
rect 539 2741 541 2748
rect 549 2741 553 2748
rect 539 2735 553 2741
rect 560 2747 579 2750
rect 560 2738 563 2747
rect 573 2738 579 2747
rect 560 2735 579 2738
rect 598 2749 617 2750
rect 598 2741 604 2749
rect 612 2741 617 2749
rect 598 2735 617 2741
rect 624 2748 638 2750
rect 764 2755 781 2759
rect 624 2740 627 2748
rect 635 2740 638 2748
rect 624 2735 638 2740
rect 661 2748 680 2749
rect 661 2740 667 2748
rect 675 2740 680 2748
rect 661 2734 680 2740
rect 687 2747 701 2749
rect 687 2739 690 2747
rect 698 2739 701 2747
rect 764 2745 766 2755
rect 776 2745 781 2755
rect 764 2743 781 2745
rect 789 2756 804 2759
rect 789 2746 791 2756
rect 801 2746 804 2756
rect 789 2743 804 2746
rect 687 2734 701 2739
rect 462 2695 464 2704
rect 470 2695 472 2704
rect 480 2695 485 2704
rect 519 2589 533 2591
rect 519 2582 521 2589
rect 529 2582 533 2589
rect 519 2576 533 2582
rect 540 2588 559 2591
rect 540 2579 543 2588
rect 553 2579 559 2588
rect 540 2576 559 2579
rect 578 2590 597 2591
rect 578 2582 584 2590
rect 592 2582 597 2590
rect 578 2576 597 2582
rect 604 2589 618 2591
rect 604 2581 607 2589
rect 615 2581 618 2589
rect 604 2576 618 2581
rect 641 2589 660 2590
rect 641 2581 647 2589
rect 655 2581 660 2589
rect 641 2575 660 2581
rect 667 2588 681 2590
rect 784 2594 801 2598
rect 667 2580 670 2588
rect 678 2580 681 2588
rect 667 2575 681 2580
rect 709 2587 728 2588
rect 709 2579 715 2587
rect 723 2579 728 2587
rect 709 2573 728 2579
rect 735 2586 749 2588
rect 735 2578 738 2586
rect 746 2578 749 2586
rect 784 2584 786 2594
rect 796 2584 801 2594
rect 784 2582 801 2584
rect 809 2595 824 2598
rect 809 2585 811 2595
rect 821 2585 824 2595
rect 809 2582 824 2585
rect 735 2573 749 2578
rect 461 2540 463 2549
rect 469 2540 471 2549
rect 479 2540 484 2549
rect 528 2370 542 2372
rect 528 2363 530 2370
rect 538 2363 542 2370
rect 528 2357 542 2363
rect 549 2369 568 2372
rect 549 2360 552 2369
rect 562 2360 568 2369
rect 549 2357 568 2360
rect 587 2371 606 2372
rect 587 2363 593 2371
rect 601 2363 606 2371
rect 587 2357 606 2363
rect 613 2370 627 2372
rect 613 2362 616 2370
rect 624 2362 627 2370
rect 613 2357 627 2362
rect 650 2370 669 2371
rect 650 2362 656 2370
rect 664 2362 669 2370
rect 650 2356 669 2362
rect 676 2369 690 2371
rect 676 2361 679 2369
rect 687 2361 690 2369
rect 676 2356 690 2361
rect 718 2368 737 2369
rect 718 2360 724 2368
rect 732 2360 737 2368
rect 718 2354 737 2360
rect 744 2367 758 2369
rect 854 2374 871 2378
rect 744 2359 747 2367
rect 755 2359 758 2367
rect 744 2354 758 2359
rect 777 2367 796 2368
rect 777 2359 783 2367
rect 791 2359 796 2367
rect 777 2353 796 2359
rect 803 2366 817 2368
rect 803 2358 806 2366
rect 814 2358 817 2366
rect 854 2364 856 2374
rect 866 2364 871 2374
rect 854 2362 871 2364
rect 879 2375 894 2378
rect 879 2365 881 2375
rect 891 2365 894 2375
rect 879 2362 894 2365
rect 803 2353 817 2358
rect 461 2308 463 2317
rect 469 2308 471 2317
rect 479 2308 484 2317
rect 1146 1990 1148 1999
rect 1154 1990 1156 1999
rect 1164 1990 1169 1999
rect 408 1980 422 1982
rect 408 1973 410 1980
rect 418 1973 422 1980
rect 408 1967 422 1973
rect 429 1979 448 1982
rect 429 1970 432 1979
rect 442 1970 448 1979
rect 429 1967 448 1970
rect 467 1981 486 1982
rect 467 1973 473 1981
rect 481 1973 486 1981
rect 467 1967 486 1973
rect 493 1980 507 1982
rect 493 1972 496 1980
rect 504 1972 507 1980
rect 493 1967 507 1972
rect 611 1980 625 1982
rect 611 1973 613 1980
rect 621 1973 625 1980
rect 611 1967 625 1973
rect 632 1979 651 1982
rect 632 1970 635 1979
rect 645 1970 651 1979
rect 632 1967 651 1970
rect 670 1981 689 1982
rect 670 1973 676 1981
rect 684 1973 689 1981
rect 670 1967 689 1973
rect 696 1980 710 1982
rect 696 1972 699 1980
rect 707 1972 710 1980
rect 696 1967 710 1972
rect 798 1980 812 1982
rect 798 1973 800 1980
rect 808 1973 812 1980
rect 798 1967 812 1973
rect 819 1979 838 1982
rect 819 1970 822 1979
rect 832 1970 838 1979
rect 819 1967 838 1970
rect 857 1981 876 1982
rect 857 1973 863 1981
rect 871 1973 876 1981
rect 857 1967 876 1973
rect 883 1980 897 1982
rect 883 1972 886 1980
rect 894 1972 897 1980
rect 883 1967 897 1972
rect 979 1980 993 1982
rect 979 1973 981 1980
rect 989 1973 993 1980
rect 979 1967 993 1973
rect 1000 1979 1019 1982
rect 1000 1970 1003 1979
rect 1013 1970 1019 1979
rect 1000 1967 1019 1970
rect 1038 1981 1057 1982
rect 1038 1973 1044 1981
rect 1052 1973 1057 1981
rect 1038 1967 1057 1973
rect 1064 1980 1078 1982
rect 1064 1972 1067 1980
rect 1075 1972 1078 1980
rect 1064 1967 1078 1972
rect 1148 1698 1150 1707
rect 1156 1698 1158 1707
rect 1166 1698 1171 1707
rect 414 1691 428 1693
rect 414 1684 416 1691
rect 424 1684 428 1691
rect 414 1678 428 1684
rect 435 1690 454 1693
rect 435 1681 438 1690
rect 448 1681 454 1690
rect 435 1678 454 1681
rect 473 1692 492 1693
rect 473 1684 479 1692
rect 487 1684 492 1692
rect 473 1678 492 1684
rect 499 1691 513 1693
rect 499 1683 502 1691
rect 510 1683 513 1691
rect 499 1678 513 1683
rect 617 1691 631 1693
rect 617 1684 619 1691
rect 627 1684 631 1691
rect 617 1678 631 1684
rect 638 1690 657 1693
rect 638 1681 641 1690
rect 651 1681 657 1690
rect 638 1678 657 1681
rect 676 1692 695 1693
rect 676 1684 682 1692
rect 690 1684 695 1692
rect 676 1678 695 1684
rect 702 1691 716 1693
rect 702 1683 705 1691
rect 713 1683 716 1691
rect 702 1678 716 1683
rect 804 1691 818 1693
rect 804 1684 806 1691
rect 814 1684 818 1691
rect 804 1678 818 1684
rect 825 1690 844 1693
rect 825 1681 828 1690
rect 838 1681 844 1690
rect 825 1678 844 1681
rect 863 1692 882 1693
rect 863 1684 869 1692
rect 877 1684 882 1692
rect 863 1678 882 1684
rect 889 1691 903 1693
rect 889 1683 892 1691
rect 900 1683 903 1691
rect 889 1678 903 1683
rect 985 1691 999 1693
rect 985 1684 987 1691
rect 995 1684 999 1691
rect 985 1678 999 1684
rect 1006 1690 1025 1693
rect 1006 1681 1009 1690
rect 1019 1681 1025 1690
rect 1006 1678 1025 1681
rect 1044 1692 1063 1693
rect 1044 1684 1050 1692
rect 1058 1684 1063 1692
rect 1044 1678 1063 1684
rect 1070 1691 1084 1693
rect 1070 1683 1073 1691
rect 1081 1683 1084 1691
rect 1070 1678 1084 1683
rect 1173 1381 1175 1390
rect 1181 1381 1183 1390
rect 1191 1381 1196 1390
rect 434 1374 448 1376
rect 434 1367 436 1374
rect 444 1367 448 1374
rect 434 1361 448 1367
rect 455 1373 474 1376
rect 455 1364 458 1373
rect 468 1364 474 1373
rect 455 1361 474 1364
rect 493 1375 512 1376
rect 493 1367 499 1375
rect 507 1367 512 1375
rect 493 1361 512 1367
rect 519 1374 533 1376
rect 519 1366 522 1374
rect 530 1366 533 1374
rect 519 1361 533 1366
rect 637 1374 651 1376
rect 637 1367 639 1374
rect 647 1367 651 1374
rect 637 1361 651 1367
rect 658 1373 677 1376
rect 658 1364 661 1373
rect 671 1364 677 1373
rect 658 1361 677 1364
rect 696 1375 715 1376
rect 696 1367 702 1375
rect 710 1367 715 1375
rect 696 1361 715 1367
rect 722 1374 736 1376
rect 722 1366 725 1374
rect 733 1366 736 1374
rect 722 1361 736 1366
rect 824 1374 838 1376
rect 824 1367 826 1374
rect 834 1367 838 1374
rect 824 1361 838 1367
rect 845 1373 864 1376
rect 845 1364 848 1373
rect 858 1364 864 1373
rect 845 1361 864 1364
rect 883 1375 902 1376
rect 883 1367 889 1375
rect 897 1367 902 1375
rect 883 1361 902 1367
rect 909 1374 923 1376
rect 909 1366 912 1374
rect 920 1366 923 1374
rect 909 1361 923 1366
rect 1005 1374 1019 1376
rect 1005 1367 1007 1374
rect 1015 1367 1019 1374
rect 1005 1361 1019 1367
rect 1026 1373 1045 1376
rect 1026 1364 1029 1373
rect 1039 1364 1045 1373
rect 1026 1361 1045 1364
rect 1064 1375 1083 1376
rect 1064 1367 1070 1375
rect 1078 1367 1083 1375
rect 1064 1361 1083 1367
rect 1090 1374 1104 1376
rect 1090 1366 1093 1374
rect 1101 1366 1104 1374
rect 1090 1361 1104 1366
rect 1182 1090 1184 1099
rect 1190 1090 1192 1099
rect 1200 1090 1205 1099
rect 432 1083 446 1085
rect 432 1076 434 1083
rect 442 1076 446 1083
rect 432 1070 446 1076
rect 453 1082 472 1085
rect 453 1073 456 1082
rect 466 1073 472 1082
rect 453 1070 472 1073
rect 491 1084 510 1085
rect 491 1076 497 1084
rect 505 1076 510 1084
rect 491 1070 510 1076
rect 517 1083 531 1085
rect 517 1075 520 1083
rect 528 1075 531 1083
rect 517 1070 531 1075
rect 635 1083 649 1085
rect 635 1076 637 1083
rect 645 1076 649 1083
rect 635 1070 649 1076
rect 656 1082 675 1085
rect 656 1073 659 1082
rect 669 1073 675 1082
rect 656 1070 675 1073
rect 694 1084 713 1085
rect 694 1076 700 1084
rect 708 1076 713 1084
rect 694 1070 713 1076
rect 720 1083 734 1085
rect 720 1075 723 1083
rect 731 1075 734 1083
rect 720 1070 734 1075
rect 822 1083 836 1085
rect 822 1076 824 1083
rect 832 1076 836 1083
rect 822 1070 836 1076
rect 843 1082 862 1085
rect 843 1073 846 1082
rect 856 1073 862 1082
rect 843 1070 862 1073
rect 881 1084 900 1085
rect 881 1076 887 1084
rect 895 1076 900 1084
rect 881 1070 900 1076
rect 907 1083 921 1085
rect 907 1075 910 1083
rect 918 1075 921 1083
rect 907 1070 921 1075
rect 1003 1083 1017 1085
rect 1003 1076 1005 1083
rect 1013 1076 1017 1083
rect 1003 1070 1017 1076
rect 1024 1082 1043 1085
rect 1024 1073 1027 1082
rect 1037 1073 1043 1082
rect 1024 1070 1043 1073
rect 1062 1084 1081 1085
rect 1062 1076 1068 1084
rect 1076 1076 1081 1084
rect 1062 1070 1081 1076
rect 1088 1083 1102 1085
rect 1088 1075 1091 1083
rect 1099 1075 1102 1083
rect 1088 1070 1102 1075
rect 485 651 499 653
rect 485 644 487 651
rect 495 644 499 651
rect 485 638 499 644
rect 506 650 525 653
rect 506 641 509 650
rect 519 641 525 650
rect 506 638 525 641
rect 544 652 563 653
rect 544 644 550 652
rect 558 644 563 652
rect 544 638 563 644
rect 570 651 584 653
rect 570 643 573 651
rect 581 643 584 651
rect 570 638 584 643
rect 655 644 672 648
rect 655 634 657 644
rect 667 634 672 644
rect 655 632 672 634
rect 680 645 695 648
rect 680 635 682 645
rect 692 635 695 645
rect 680 632 695 635
rect 406 591 408 600
rect 414 591 416 600
rect 424 591 429 600
rect 485 482 499 484
rect 485 475 487 482
rect 495 475 499 482
rect 485 469 499 475
rect 506 481 525 484
rect 506 472 509 481
rect 519 472 525 481
rect 506 469 525 472
rect 544 483 563 484
rect 544 475 550 483
rect 558 475 563 483
rect 544 469 563 475
rect 570 482 584 484
rect 710 489 727 493
rect 570 474 573 482
rect 581 474 584 482
rect 570 469 584 474
rect 607 482 626 483
rect 607 474 613 482
rect 621 474 626 482
rect 607 468 626 474
rect 633 481 647 483
rect 633 473 636 481
rect 644 473 647 481
rect 710 479 712 489
rect 722 479 727 489
rect 710 477 727 479
rect 735 490 750 493
rect 735 480 737 490
rect 747 480 750 490
rect 735 477 750 480
rect 633 468 647 473
rect 2288 2729 2290 2738
rect 2296 2729 2298 2738
rect 2306 2729 2311 2738
rect 2078 2708 2092 2710
rect 2078 2701 2080 2708
rect 2088 2701 2092 2708
rect 2078 2695 2092 2701
rect 2099 2707 2118 2710
rect 2099 2698 2102 2707
rect 2112 2698 2118 2707
rect 2099 2695 2118 2698
rect 2137 2709 2156 2710
rect 2137 2701 2143 2709
rect 2151 2701 2156 2709
rect 2137 2695 2156 2701
rect 2164 2708 2177 2710
rect 2164 2700 2166 2708
rect 2174 2700 2177 2708
rect 2164 2695 2177 2700
rect 2213 2709 2229 2711
rect 2213 2701 2219 2709
rect 2227 2701 2229 2709
rect 2213 2696 2229 2701
rect 2237 2708 2255 2711
rect 2237 2699 2239 2708
rect 2249 2699 2255 2708
rect 2237 2696 2255 2699
rect 1635 1417 1637 1426
rect 1643 1417 1645 1426
rect 1653 1417 1658 1426
rect 2288 1430 2290 1439
rect 2296 1430 2298 1439
rect 2306 1430 2311 1439
rect 2078 1409 2092 1411
rect 1357 1406 1371 1408
rect 1357 1399 1359 1406
rect 1367 1399 1371 1406
rect 1357 1393 1371 1399
rect 1378 1405 1397 1408
rect 1378 1396 1381 1405
rect 1391 1396 1397 1405
rect 1378 1393 1397 1396
rect 1416 1407 1435 1408
rect 1416 1399 1422 1407
rect 1430 1399 1435 1407
rect 1416 1393 1435 1399
rect 1442 1406 1456 1408
rect 1442 1398 1445 1406
rect 1453 1398 1456 1406
rect 1442 1393 1456 1398
rect 1492 1407 1508 1409
rect 1492 1399 1498 1407
rect 1506 1399 1508 1407
rect 1492 1394 1508 1399
rect 1515 1406 1534 1409
rect 1515 1397 1518 1406
rect 1528 1397 1534 1406
rect 1515 1394 1534 1397
rect 1553 1408 1572 1409
rect 1553 1400 1559 1408
rect 1567 1400 1572 1408
rect 1553 1394 1572 1400
rect 1579 1407 1593 1409
rect 1579 1399 1582 1407
rect 1590 1399 1593 1407
rect 1579 1394 1593 1399
rect 2078 1402 2080 1409
rect 2088 1402 2092 1409
rect 2078 1396 2092 1402
rect 2099 1408 2118 1411
rect 2099 1399 2102 1408
rect 2112 1399 2118 1408
rect 2099 1396 2118 1399
rect 2137 1410 2156 1411
rect 2137 1402 2143 1410
rect 2151 1402 2156 1410
rect 2137 1396 2156 1402
rect 2163 1409 2177 1411
rect 2163 1401 2166 1409
rect 2174 1401 2177 1409
rect 2163 1396 2177 1401
rect 2213 1410 2229 1412
rect 2213 1402 2219 1410
rect 2227 1402 2229 1410
rect 2213 1397 2229 1402
rect 2236 1409 2255 1412
rect 2236 1400 2239 1409
rect 2249 1400 2255 1409
rect 2236 1397 2255 1400
rect 408 429 410 438
rect 416 429 418 438
rect 426 429 431 438
rect 465 323 479 325
rect 465 316 467 323
rect 475 316 479 323
rect 465 310 479 316
rect 486 322 505 325
rect 486 313 489 322
rect 499 313 505 322
rect 486 310 505 313
rect 524 324 543 325
rect 524 316 530 324
rect 538 316 543 324
rect 524 310 543 316
rect 550 323 564 325
rect 550 315 553 323
rect 561 315 564 323
rect 550 310 564 315
rect 587 323 606 324
rect 587 315 593 323
rect 601 315 606 323
rect 587 309 606 315
rect 613 322 627 324
rect 730 328 747 332
rect 613 314 616 322
rect 624 314 627 322
rect 613 309 627 314
rect 655 321 674 322
rect 655 313 661 321
rect 669 313 674 321
rect 655 307 674 313
rect 681 320 695 322
rect 681 312 684 320
rect 692 312 695 320
rect 730 318 732 328
rect 742 318 747 328
rect 730 316 747 318
rect 755 329 770 332
rect 755 319 757 329
rect 767 319 770 329
rect 755 316 770 319
rect 681 307 695 312
rect 407 274 409 283
rect 415 274 417 283
rect 425 274 430 283
rect 474 104 488 106
rect 474 97 476 104
rect 484 97 488 104
rect 474 91 488 97
rect 495 103 514 106
rect 495 94 498 103
rect 508 94 514 103
rect 495 91 514 94
rect 533 105 552 106
rect 533 97 539 105
rect 547 97 552 105
rect 533 91 552 97
rect 559 104 573 106
rect 559 96 562 104
rect 570 96 573 104
rect 559 91 573 96
rect 596 104 615 105
rect 596 96 602 104
rect 610 96 615 104
rect 596 90 615 96
rect 622 103 636 105
rect 622 95 625 103
rect 633 95 636 103
rect 622 90 636 95
rect 664 102 683 103
rect 664 94 670 102
rect 678 94 683 102
rect 664 88 683 94
rect 690 101 704 103
rect 800 108 817 112
rect 690 93 693 101
rect 701 93 704 101
rect 690 88 704 93
rect 723 101 742 102
rect 723 93 729 101
rect 737 93 742 101
rect 723 87 742 93
rect 749 100 763 102
rect 749 92 752 100
rect 760 92 763 100
rect 800 98 802 108
rect 812 98 817 108
rect 800 96 817 98
rect 825 109 840 112
rect 825 99 827 109
rect 837 99 840 109
rect 825 96 840 99
rect 749 87 763 92
rect 5045 971 5056 974
rect 5045 966 5047 971
rect 5053 966 5056 971
rect 5045 963 5056 966
rect 5062 972 5078 974
rect 5062 966 5066 972
rect 5073 966 5078 972
rect 5062 963 5078 966
rect 5083 971 5097 974
rect 5083 966 5087 971
rect 5093 966 5097 971
rect 5083 963 5097 966
rect 5103 973 5114 974
rect 5103 966 5104 973
rect 5111 966 5114 973
rect 5103 963 5114 966
rect 5124 971 5138 974
rect 5124 965 5128 971
rect 5134 965 5138 971
rect 5124 963 5138 965
rect 5144 972 5157 974
rect 5144 966 5146 972
rect 5153 966 5157 972
rect 5144 963 5157 966
rect 5164 971 5180 974
rect 5164 966 5170 971
rect 5176 966 5180 971
rect 5164 963 5180 966
rect 5186 972 5197 974
rect 5186 966 5188 972
rect 5195 966 5197 972
rect 5186 963 5197 966
rect 4788 934 4799 937
rect 4788 929 4790 934
rect 4796 929 4799 934
rect 4788 926 4799 929
rect 4805 935 4821 937
rect 4805 929 4809 935
rect 4816 929 4821 935
rect 4805 926 4821 929
rect 4826 934 4840 937
rect 4826 929 4830 934
rect 4836 929 4840 934
rect 4826 926 4840 929
rect 4846 936 4857 937
rect 4846 929 4847 936
rect 4854 929 4857 936
rect 4846 926 4857 929
rect 4867 934 4881 937
rect 4867 928 4871 934
rect 4877 928 4881 934
rect 4867 926 4881 928
rect 4887 935 4900 937
rect 4887 929 4889 935
rect 4896 929 4900 935
rect 4887 926 4900 929
rect 4907 934 4923 937
rect 4907 929 4913 934
rect 4919 929 4923 934
rect 4907 926 4923 929
rect 4929 935 4940 937
rect 4929 929 4931 935
rect 4938 929 4940 935
rect 4929 926 4940 929
rect 4544 779 4555 782
rect 4544 774 4546 779
rect 4552 774 4555 779
rect 4544 771 4555 774
rect 4561 780 4577 782
rect 4561 774 4565 780
rect 4572 774 4577 780
rect 4561 771 4577 774
rect 4582 779 4596 782
rect 4582 774 4586 779
rect 4592 774 4596 779
rect 4582 771 4596 774
rect 4602 781 4613 782
rect 4602 774 4603 781
rect 4610 774 4613 781
rect 4602 771 4613 774
rect 4623 779 4637 782
rect 4623 773 4627 779
rect 4633 773 4637 779
rect 4623 771 4637 773
rect 4643 780 4656 782
rect 4643 774 4645 780
rect 4652 774 4656 780
rect 4643 771 4656 774
rect 4663 779 4679 782
rect 4663 774 4669 779
rect 4675 774 4679 779
rect 4663 771 4679 774
rect 4685 780 4696 782
rect 4685 774 4687 780
rect 4694 774 4696 780
rect 4685 771 4696 774
rect 1565 585 1576 588
rect 1565 580 1567 585
rect 1573 580 1576 585
rect 1565 577 1576 580
rect 1582 586 1598 588
rect 1582 580 1586 586
rect 1593 580 1598 586
rect 1582 577 1598 580
rect 1603 585 1617 588
rect 1603 580 1607 585
rect 1613 580 1617 585
rect 1603 577 1617 580
rect 1623 586 1636 588
rect 1623 580 1626 586
rect 1633 580 1636 586
rect 1623 577 1636 580
rect 1642 585 1656 588
rect 1642 579 1646 585
rect 1652 579 1656 585
rect 1642 577 1656 579
rect 1662 587 1675 588
rect 1662 580 1665 587
rect 1672 580 1675 587
rect 1662 577 1675 580
rect 1685 585 1699 588
rect 1685 579 1689 585
rect 1695 579 1699 585
rect 1685 577 1699 579
rect 1705 586 1718 588
rect 1705 580 1707 586
rect 1714 580 1718 586
rect 1705 577 1718 580
rect 1725 585 1741 588
rect 1725 580 1731 585
rect 1737 580 1741 585
rect 1725 577 1741 580
rect 1747 586 1758 588
rect 1747 580 1749 586
rect 1756 580 1758 586
rect 2288 599 2290 608
rect 2296 599 2298 608
rect 2306 599 2311 608
rect 1747 577 1758 580
rect 2078 578 2092 580
rect 407 42 409 51
rect 415 42 417 51
rect 425 42 430 51
rect 2078 571 2080 578
rect 2088 571 2092 578
rect 2078 565 2092 571
rect 2099 577 2118 580
rect 2099 568 2102 577
rect 2112 568 2118 577
rect 2099 565 2118 568
rect 2137 579 2156 580
rect 2137 571 2143 579
rect 2151 571 2156 579
rect 2137 565 2156 571
rect 2163 578 2177 580
rect 2163 570 2166 578
rect 2174 570 2177 578
rect 2163 565 2177 570
rect 2213 579 2229 581
rect 2213 571 2219 579
rect 2227 571 2229 579
rect 2213 566 2229 571
rect 2236 578 2255 581
rect 2236 569 2239 578
rect 2249 569 2255 578
rect 2236 566 2255 569
rect 691 -396 705 -394
rect 691 -403 693 -396
rect 701 -403 705 -396
rect 691 -409 705 -403
rect 712 -397 731 -394
rect 712 -406 715 -397
rect 725 -406 731 -397
rect 712 -409 731 -406
rect 750 -395 769 -394
rect 750 -403 756 -395
rect 764 -403 769 -395
rect 750 -409 769 -403
rect 776 -396 790 -394
rect 776 -404 779 -396
rect 787 -404 790 -396
rect 776 -409 790 -404
rect 861 -403 878 -399
rect 861 -413 863 -403
rect 873 -413 878 -403
rect 861 -415 878 -413
rect 886 -402 901 -399
rect 886 -412 888 -402
rect 898 -412 901 -402
rect 886 -415 901 -412
rect 1489 -418 1491 -409
rect 1497 -418 1499 -409
rect 1507 -418 1512 -409
rect 1279 -439 1293 -437
rect 1279 -446 1281 -439
rect 1289 -446 1293 -439
rect 1279 -452 1293 -446
rect 1300 -440 1319 -437
rect 1300 -449 1303 -440
rect 1313 -449 1319 -440
rect 1300 -452 1319 -449
rect 1338 -438 1357 -437
rect 1338 -446 1344 -438
rect 1352 -446 1357 -438
rect 1338 -452 1357 -446
rect 1364 -439 1378 -437
rect 1364 -447 1367 -439
rect 1375 -447 1378 -439
rect 1364 -452 1378 -447
rect 1414 -438 1430 -436
rect 1414 -446 1420 -438
rect 1428 -446 1430 -438
rect 1414 -451 1430 -446
rect 1438 -439 1456 -436
rect 1438 -448 1440 -439
rect 1450 -448 1456 -439
rect 1438 -451 1456 -448
rect 693 -594 707 -592
rect 693 -601 695 -594
rect 703 -601 707 -594
rect 693 -607 707 -601
rect 714 -595 733 -592
rect 714 -604 717 -595
rect 727 -604 733 -595
rect 714 -607 733 -604
rect 752 -593 771 -592
rect 752 -601 758 -593
rect 766 -601 771 -593
rect 752 -607 771 -601
rect 778 -594 792 -592
rect 778 -602 781 -594
rect 789 -602 792 -594
rect 778 -607 792 -602
rect 863 -601 880 -597
rect 863 -611 865 -601
rect 875 -611 880 -601
rect 863 -613 880 -611
rect 888 -600 903 -597
rect 888 -610 890 -600
rect 900 -610 903 -600
rect 888 -613 903 -610
rect 1489 -608 1491 -599
rect 1497 -608 1499 -599
rect 1507 -608 1512 -599
rect 1279 -629 1293 -627
rect 1279 -636 1281 -629
rect 1289 -636 1293 -629
rect 1279 -642 1293 -636
rect 1300 -630 1319 -627
rect 1300 -639 1303 -630
rect 1313 -639 1319 -630
rect 1300 -642 1319 -639
rect 1338 -628 1357 -627
rect 1338 -636 1344 -628
rect 1352 -636 1357 -628
rect 1338 -642 1357 -636
rect 1364 -629 1378 -627
rect 1364 -637 1367 -629
rect 1375 -637 1378 -629
rect 1364 -642 1378 -637
rect 1414 -628 1430 -626
rect 1414 -636 1420 -628
rect 1428 -636 1430 -628
rect 1414 -641 1430 -636
rect 1437 -629 1456 -626
rect 1437 -638 1440 -629
rect 1450 -638 1456 -629
rect 1437 -641 1456 -638
rect 693 -792 707 -790
rect 693 -799 695 -792
rect 703 -799 707 -792
rect 693 -805 707 -799
rect 714 -793 733 -790
rect 714 -802 717 -793
rect 727 -802 733 -793
rect 714 -805 733 -802
rect 752 -791 771 -790
rect 752 -799 758 -791
rect 766 -799 771 -791
rect 752 -805 771 -799
rect 778 -792 792 -790
rect 778 -800 781 -792
rect 789 -800 792 -792
rect 778 -805 792 -800
rect 863 -799 880 -795
rect 863 -809 865 -799
rect 875 -809 880 -799
rect 863 -811 880 -809
rect 888 -798 903 -795
rect 888 -808 890 -798
rect 900 -808 903 -798
rect 888 -811 903 -808
rect 5246 598 5257 601
rect 5246 593 5248 598
rect 5254 593 5257 598
rect 5246 590 5257 593
rect 5263 599 5279 601
rect 5263 593 5267 599
rect 5274 593 5279 599
rect 5263 590 5279 593
rect 5284 598 5298 601
rect 5284 593 5288 598
rect 5294 593 5298 598
rect 5284 590 5298 593
rect 5304 599 5317 601
rect 5304 593 5307 599
rect 5314 593 5317 599
rect 5304 590 5317 593
rect 5333 598 5349 601
rect 5333 593 5339 598
rect 5345 593 5349 598
rect 5333 590 5349 593
rect 5355 599 5366 601
rect 5355 593 5357 599
rect 5364 593 5366 599
rect 5355 590 5366 593
rect 1489 -814 1491 -805
rect 1497 -814 1499 -805
rect 1507 -814 1512 -805
rect 1279 -835 1293 -833
rect 1279 -842 1281 -835
rect 1289 -842 1293 -835
rect 1279 -848 1293 -842
rect 1300 -836 1319 -833
rect 1300 -845 1303 -836
rect 1313 -845 1319 -836
rect 1300 -848 1319 -845
rect 1338 -834 1357 -833
rect 1338 -842 1344 -834
rect 1352 -842 1357 -834
rect 1338 -848 1357 -842
rect 1364 -835 1378 -833
rect 1364 -843 1367 -835
rect 1375 -843 1378 -835
rect 1364 -848 1378 -843
rect 1414 -834 1430 -832
rect 1414 -842 1420 -834
rect 1428 -842 1430 -834
rect 1414 -847 1430 -842
rect 1438 -835 1456 -832
rect 1438 -844 1440 -835
rect 1450 -844 1456 -835
rect 1438 -847 1456 -844
rect 693 -987 707 -985
rect 693 -994 695 -987
rect 703 -994 707 -987
rect 693 -1000 707 -994
rect 714 -988 733 -985
rect 714 -997 717 -988
rect 727 -997 733 -988
rect 714 -1000 733 -997
rect 752 -986 771 -985
rect 752 -994 758 -986
rect 766 -994 771 -986
rect 752 -1000 771 -994
rect 778 -987 792 -985
rect 778 -995 781 -987
rect 789 -995 792 -987
rect 778 -1000 792 -995
rect 863 -994 880 -990
rect 863 -1004 865 -994
rect 875 -1004 880 -994
rect 863 -1006 880 -1004
rect 888 -993 903 -990
rect 888 -1003 890 -993
rect 900 -1003 903 -993
rect 888 -1006 903 -1003
rect 1489 -1004 1491 -995
rect 1497 -1004 1499 -995
rect 1507 -1004 1512 -995
rect 1279 -1025 1293 -1023
rect 1279 -1032 1281 -1025
rect 1289 -1032 1293 -1025
rect 1279 -1038 1293 -1032
rect 1300 -1026 1319 -1023
rect 1300 -1035 1303 -1026
rect 1313 -1035 1319 -1026
rect 1300 -1038 1319 -1035
rect 1338 -1024 1357 -1023
rect 1338 -1032 1344 -1024
rect 1352 -1032 1357 -1024
rect 1338 -1038 1357 -1032
rect 1364 -1025 1378 -1023
rect 1364 -1033 1367 -1025
rect 1375 -1033 1378 -1025
rect 1364 -1038 1378 -1033
rect 1414 -1024 1430 -1022
rect 1414 -1032 1420 -1024
rect 1428 -1032 1430 -1024
rect 1414 -1037 1430 -1032
rect 1437 -1025 1456 -1022
rect 1437 -1034 1440 -1025
rect 1450 -1034 1456 -1025
rect 1437 -1037 1456 -1034
<< pdiffusion >>
rect -662 5980 -648 5982
rect -662 5974 -659 5980
rect -652 5974 -648 5980
rect -662 5967 -648 5974
rect -641 5978 -622 5982
rect -641 5970 -637 5978
rect -628 5970 -622 5978
rect -641 5967 -622 5970
rect -595 5978 -584 5982
rect -595 5971 -593 5978
rect -585 5971 -584 5978
rect -595 5967 -584 5971
rect -577 5976 -555 5982
rect -577 5970 -574 5976
rect -566 5970 -555 5976
rect -577 5967 -555 5970
rect -459 5980 -445 5982
rect -459 5974 -456 5980
rect -449 5974 -445 5980
rect -459 5967 -445 5974
rect -438 5978 -419 5982
rect -438 5970 -434 5978
rect -425 5970 -419 5978
rect -438 5967 -419 5970
rect -392 5978 -381 5982
rect -392 5971 -390 5978
rect -382 5971 -381 5978
rect -392 5967 -381 5971
rect -374 5976 -352 5982
rect -374 5970 -371 5976
rect -363 5970 -352 5976
rect -374 5967 -352 5970
rect -272 5980 -258 5982
rect -272 5974 -269 5980
rect -262 5974 -258 5980
rect -272 5967 -258 5974
rect -251 5978 -232 5982
rect -251 5970 -247 5978
rect -238 5970 -232 5978
rect -251 5967 -232 5970
rect -205 5978 -194 5982
rect -205 5971 -203 5978
rect -195 5971 -194 5978
rect -205 5967 -194 5971
rect -187 5976 -165 5982
rect -187 5970 -184 5976
rect -176 5970 -165 5976
rect -187 5967 -165 5970
rect -91 5980 -77 5982
rect -91 5974 -88 5980
rect -81 5974 -77 5980
rect -91 5967 -77 5974
rect -70 5978 -51 5982
rect -70 5970 -66 5978
rect -57 5970 -51 5978
rect -70 5967 -51 5970
rect -24 5978 -13 5982
rect -24 5971 -22 5978
rect -14 5971 -13 5978
rect -24 5967 -13 5971
rect -6 5976 16 5982
rect -6 5970 -3 5976
rect 5 5970 16 5976
rect -6 5967 16 5970
rect -634 5633 -620 5635
rect -634 5627 -631 5633
rect -624 5627 -620 5633
rect -634 5620 -620 5627
rect -613 5631 -594 5635
rect -613 5623 -609 5631
rect -600 5623 -594 5631
rect -613 5620 -594 5623
rect -567 5631 -556 5635
rect -567 5624 -565 5631
rect -557 5624 -556 5631
rect -567 5620 -556 5624
rect -549 5629 -527 5635
rect -549 5623 -546 5629
rect -538 5623 -527 5629
rect -549 5620 -527 5623
rect -431 5633 -417 5635
rect -431 5627 -428 5633
rect -421 5627 -417 5633
rect -431 5620 -417 5627
rect -410 5631 -391 5635
rect -410 5623 -406 5631
rect -397 5623 -391 5631
rect -410 5620 -391 5623
rect -364 5631 -353 5635
rect -364 5624 -362 5631
rect -354 5624 -353 5631
rect -364 5620 -353 5624
rect -346 5629 -324 5635
rect -346 5623 -343 5629
rect -335 5623 -324 5629
rect -346 5620 -324 5623
rect -244 5633 -230 5635
rect -244 5627 -241 5633
rect -234 5627 -230 5633
rect -244 5620 -230 5627
rect -223 5631 -204 5635
rect -223 5623 -219 5631
rect -210 5623 -204 5631
rect -223 5620 -204 5623
rect -177 5631 -166 5635
rect -177 5624 -175 5631
rect -167 5624 -166 5631
rect -177 5620 -166 5624
rect -159 5629 -137 5635
rect -159 5623 -156 5629
rect -148 5623 -137 5629
rect -159 5620 -137 5623
rect -63 5633 -49 5635
rect -63 5627 -60 5633
rect -53 5627 -49 5633
rect -63 5620 -49 5627
rect -42 5631 -23 5635
rect -42 5623 -38 5631
rect -29 5623 -23 5631
rect -42 5620 -23 5623
rect 4 5631 15 5635
rect 4 5624 6 5631
rect 14 5624 15 5631
rect 4 5620 15 5624
rect 22 5629 44 5635
rect 22 5623 25 5629
rect 33 5623 44 5629
rect 22 5620 44 5623
rect -634 5247 -620 5249
rect -634 5241 -631 5247
rect -624 5241 -620 5247
rect -634 5234 -620 5241
rect -613 5245 -594 5249
rect -613 5237 -609 5245
rect -600 5237 -594 5245
rect -613 5234 -594 5237
rect -567 5245 -556 5249
rect -567 5238 -565 5245
rect -557 5238 -556 5245
rect -567 5234 -556 5238
rect -549 5243 -527 5249
rect -549 5237 -546 5243
rect -538 5237 -527 5243
rect -549 5234 -527 5237
rect -431 5247 -417 5249
rect -431 5241 -428 5247
rect -421 5241 -417 5247
rect -431 5234 -417 5241
rect -410 5245 -391 5249
rect -410 5237 -406 5245
rect -397 5237 -391 5245
rect -410 5234 -391 5237
rect -364 5245 -353 5249
rect -364 5238 -362 5245
rect -354 5238 -353 5245
rect -364 5234 -353 5238
rect -346 5243 -324 5249
rect -346 5237 -343 5243
rect -335 5237 -324 5243
rect -346 5234 -324 5237
rect -244 5247 -230 5249
rect -244 5241 -241 5247
rect -234 5241 -230 5247
rect -244 5234 -230 5241
rect -223 5245 -204 5249
rect -223 5237 -219 5245
rect -210 5237 -204 5245
rect -223 5234 -204 5237
rect -177 5245 -166 5249
rect -177 5238 -175 5245
rect -167 5238 -166 5245
rect -177 5234 -166 5238
rect -159 5243 -137 5249
rect -159 5237 -156 5243
rect -148 5237 -137 5243
rect -159 5234 -137 5237
rect -63 5247 -49 5249
rect -63 5241 -60 5247
rect -53 5241 -49 5247
rect -63 5234 -49 5241
rect -42 5245 -23 5249
rect -42 5237 -38 5245
rect -29 5237 -23 5245
rect -42 5234 -23 5237
rect 4 5245 15 5249
rect 4 5238 6 5245
rect 14 5238 15 5245
rect 4 5234 15 5238
rect 22 5243 44 5249
rect 22 5237 25 5243
rect 33 5237 44 5243
rect 22 5234 44 5237
rect -634 4823 -620 4825
rect -634 4817 -631 4823
rect -624 4817 -620 4823
rect -634 4810 -620 4817
rect -613 4821 -594 4825
rect -613 4813 -609 4821
rect -600 4813 -594 4821
rect -613 4810 -594 4813
rect -567 4821 -556 4825
rect -567 4814 -565 4821
rect -557 4814 -556 4821
rect -567 4810 -556 4814
rect -549 4819 -527 4825
rect -549 4813 -546 4819
rect -538 4813 -527 4819
rect -549 4810 -527 4813
rect -431 4823 -417 4825
rect -431 4817 -428 4823
rect -421 4817 -417 4823
rect -431 4810 -417 4817
rect -410 4821 -391 4825
rect -410 4813 -406 4821
rect -397 4813 -391 4821
rect -410 4810 -391 4813
rect -364 4821 -353 4825
rect -364 4814 -362 4821
rect -354 4814 -353 4821
rect -364 4810 -353 4814
rect -346 4819 -324 4825
rect -346 4813 -343 4819
rect -335 4813 -324 4819
rect -346 4810 -324 4813
rect -244 4823 -230 4825
rect -244 4817 -241 4823
rect -234 4817 -230 4823
rect -244 4810 -230 4817
rect -223 4821 -204 4825
rect -223 4813 -219 4821
rect -210 4813 -204 4821
rect -223 4810 -204 4813
rect -177 4821 -166 4825
rect -177 4814 -175 4821
rect -167 4814 -166 4821
rect -177 4810 -166 4814
rect -159 4819 -137 4825
rect -159 4813 -156 4819
rect -148 4813 -137 4819
rect -159 4810 -137 4813
rect -63 4823 -49 4825
rect -63 4817 -60 4823
rect -53 4817 -49 4823
rect -63 4810 -49 4817
rect -42 4821 -23 4825
rect -42 4813 -38 4821
rect -29 4813 -23 4821
rect -42 4810 -23 4813
rect 4 4821 15 4825
rect 4 4814 6 4821
rect 14 4814 15 4821
rect 4 4810 15 4814
rect 22 4819 44 4825
rect 22 4813 25 4819
rect 33 4813 44 4819
rect 22 4810 44 4813
rect 432 5701 446 5703
rect 432 5695 435 5701
rect 442 5695 446 5701
rect 432 5688 446 5695
rect 453 5699 472 5703
rect 453 5691 457 5699
rect 466 5691 472 5699
rect 453 5688 472 5691
rect 499 5699 510 5703
rect 499 5692 501 5699
rect 509 5692 510 5699
rect 499 5688 510 5692
rect 517 5697 539 5703
rect 517 5691 520 5697
rect 528 5691 539 5697
rect 517 5688 539 5691
rect 635 5701 649 5703
rect 635 5695 638 5701
rect 645 5695 649 5701
rect 635 5688 649 5695
rect 656 5699 675 5703
rect 656 5691 660 5699
rect 669 5691 675 5699
rect 656 5688 675 5691
rect 702 5699 713 5703
rect 702 5692 704 5699
rect 712 5692 713 5699
rect 702 5688 713 5692
rect 720 5697 742 5703
rect 720 5691 723 5697
rect 731 5691 742 5697
rect 720 5688 742 5691
rect 822 5701 836 5703
rect 822 5695 825 5701
rect 832 5695 836 5701
rect 822 5688 836 5695
rect 843 5699 862 5703
rect 843 5691 847 5699
rect 856 5691 862 5699
rect 843 5688 862 5691
rect 889 5699 900 5703
rect 889 5692 891 5699
rect 899 5692 900 5699
rect 889 5688 900 5692
rect 907 5697 929 5703
rect 907 5691 910 5697
rect 918 5691 929 5697
rect 907 5688 929 5691
rect 1003 5701 1017 5703
rect 1003 5695 1006 5701
rect 1013 5695 1017 5701
rect 1003 5688 1017 5695
rect 1024 5699 1043 5703
rect 1024 5691 1028 5699
rect 1037 5691 1043 5699
rect 1024 5688 1043 5691
rect 1070 5699 1081 5703
rect 1070 5692 1072 5699
rect 1080 5692 1081 5699
rect 1070 5688 1081 5692
rect 1088 5697 1110 5703
rect 1088 5691 1091 5697
rect 1099 5691 1110 5697
rect 1088 5688 1110 5691
rect 1172 5695 1186 5697
rect 1172 5689 1175 5695
rect 1182 5689 1186 5695
rect 1172 5682 1186 5689
rect 1193 5693 1212 5697
rect 1193 5685 1197 5693
rect 1206 5685 1212 5693
rect 1193 5682 1212 5685
rect 1239 5693 1250 5697
rect 1239 5686 1241 5693
rect 1249 5686 1250 5693
rect 1239 5682 1250 5686
rect 1257 5691 1279 5697
rect 1257 5685 1260 5691
rect 1268 5685 1279 5691
rect 1257 5682 1279 5685
rect 1375 5695 1389 5697
rect 1375 5689 1378 5695
rect 1385 5689 1389 5695
rect 1375 5682 1389 5689
rect 1396 5693 1415 5697
rect 1396 5685 1400 5693
rect 1409 5685 1415 5693
rect 1396 5682 1415 5685
rect 1442 5693 1453 5697
rect 1442 5686 1444 5693
rect 1452 5686 1453 5693
rect 1442 5682 1453 5686
rect 1460 5691 1482 5697
rect 1460 5685 1463 5691
rect 1471 5685 1482 5691
rect 1460 5682 1482 5685
rect 1562 5695 1576 5697
rect 1562 5689 1565 5695
rect 1572 5689 1576 5695
rect 1562 5682 1576 5689
rect 1583 5693 1602 5697
rect 1583 5685 1587 5693
rect 1596 5685 1602 5693
rect 1583 5682 1602 5685
rect 1629 5693 1640 5697
rect 1629 5686 1631 5693
rect 1639 5686 1640 5693
rect 1629 5682 1640 5686
rect 1647 5691 1669 5697
rect 1647 5685 1650 5691
rect 1658 5685 1669 5691
rect 1647 5682 1669 5685
rect 1743 5695 1757 5697
rect 1743 5689 1746 5695
rect 1753 5689 1757 5695
rect 1743 5682 1757 5689
rect 1764 5693 1783 5697
rect 1764 5685 1768 5693
rect 1777 5685 1783 5693
rect 1764 5682 1783 5685
rect 1810 5693 1821 5697
rect 1810 5686 1812 5693
rect 1820 5686 1821 5693
rect 1810 5682 1821 5686
rect 1828 5691 1850 5697
rect 1828 5685 1831 5691
rect 1839 5685 1850 5691
rect 1828 5682 1850 5685
rect 2188 5693 2202 5695
rect 2188 5687 2191 5693
rect 2198 5687 2202 5693
rect 2188 5680 2202 5687
rect 2209 5691 2228 5695
rect 2209 5683 2213 5691
rect 2222 5683 2228 5691
rect 2209 5680 2228 5683
rect 2255 5691 2266 5695
rect 2255 5684 2257 5691
rect 2265 5684 2266 5691
rect 2255 5680 2266 5684
rect 2273 5689 2295 5695
rect 2273 5683 2276 5689
rect 2284 5683 2295 5689
rect 2273 5680 2295 5683
rect 2359 5673 2361 5683
rect 2371 5673 2375 5683
rect 2359 5667 2375 5673
rect 2383 5680 2399 5683
rect 2383 5670 2385 5680
rect 2395 5670 2399 5680
rect 2383 5667 2399 5670
rect 3040 5695 3042 5704
rect 3048 5695 3050 5704
rect 3059 5695 3063 5704
rect 3311 5618 3313 5627
rect 3319 5618 3321 5627
rect 3330 5618 3334 5627
rect 332 5409 346 5411
rect 332 5403 335 5409
rect 342 5403 346 5409
rect 332 5396 346 5403
rect 353 5407 372 5411
rect 353 5399 357 5407
rect 366 5399 372 5407
rect 353 5396 372 5399
rect 399 5407 410 5411
rect 399 5400 401 5407
rect 409 5400 410 5407
rect 399 5396 410 5400
rect 418 5405 439 5411
rect 418 5399 420 5405
rect 428 5399 439 5405
rect 418 5396 439 5399
rect 503 5389 505 5399
rect 515 5389 519 5399
rect 503 5383 519 5389
rect 527 5396 543 5399
rect 527 5386 529 5396
rect 539 5386 543 5396
rect 527 5383 543 5386
rect 615 5405 629 5407
rect 615 5399 618 5405
rect 625 5399 629 5405
rect 615 5392 629 5399
rect 636 5403 655 5407
rect 636 5395 640 5403
rect 649 5395 655 5403
rect 636 5392 655 5395
rect 682 5403 693 5407
rect 682 5396 684 5403
rect 692 5396 693 5403
rect 682 5392 693 5396
rect 700 5401 722 5407
rect 700 5395 703 5401
rect 711 5395 722 5401
rect 878 5397 889 5399
rect 700 5392 722 5395
rect 786 5385 788 5395
rect 798 5385 802 5395
rect 786 5379 802 5385
rect 810 5392 826 5395
rect 810 5382 812 5392
rect 822 5382 826 5392
rect 878 5391 880 5397
rect 886 5391 889 5397
rect 878 5388 889 5391
rect 895 5394 911 5399
rect 895 5388 899 5394
rect 905 5388 911 5394
rect 916 5394 930 5399
rect 916 5388 920 5394
rect 926 5388 930 5394
rect 936 5394 949 5399
rect 936 5388 940 5394
rect 946 5388 949 5394
rect 968 5397 981 5399
rect 968 5391 971 5397
rect 977 5391 981 5397
rect 968 5388 981 5391
rect 987 5395 1001 5399
rect 987 5389 989 5395
rect 996 5389 1001 5395
rect 987 5388 1001 5389
rect 810 5379 826 5382
rect 489 4977 503 4979
rect 489 4971 492 4977
rect 499 4971 503 4977
rect 489 4964 503 4971
rect 510 4975 529 4979
rect 510 4967 514 4975
rect 523 4967 529 4975
rect 510 4964 529 4967
rect 556 4975 567 4979
rect 556 4968 558 4975
rect 566 4968 567 4975
rect 556 4964 567 4968
rect 574 4973 596 4979
rect 574 4967 577 4973
rect 585 4967 596 4973
rect 574 4964 596 4967
rect 692 4977 706 4979
rect 692 4971 695 4977
rect 702 4971 706 4977
rect 692 4964 706 4971
rect 713 4975 732 4979
rect 713 4967 717 4975
rect 726 4967 732 4975
rect 713 4964 732 4967
rect 759 4975 770 4979
rect 759 4968 761 4975
rect 769 4968 770 4975
rect 759 4964 770 4968
rect 777 4973 799 4979
rect 777 4967 780 4973
rect 788 4967 799 4973
rect 777 4964 799 4967
rect 879 4977 893 4979
rect 879 4971 882 4977
rect 889 4971 893 4977
rect 879 4964 893 4971
rect 900 4975 919 4979
rect 900 4967 904 4975
rect 913 4967 919 4975
rect 900 4964 919 4967
rect 946 4975 957 4979
rect 946 4968 948 4975
rect 956 4968 957 4975
rect 946 4964 957 4968
rect 964 4973 986 4979
rect 964 4967 967 4973
rect 975 4967 986 4973
rect 964 4964 986 4967
rect 1060 4977 1074 4979
rect 1060 4971 1063 4977
rect 1070 4971 1074 4977
rect 1060 4964 1074 4971
rect 1081 4975 1100 4979
rect 1081 4967 1085 4975
rect 1094 4967 1100 4975
rect 1081 4964 1100 4967
rect 1127 4975 1138 4979
rect 1127 4968 1129 4975
rect 1137 4968 1138 4975
rect 1127 4964 1138 4968
rect 1145 4973 1167 4979
rect 1145 4967 1148 4973
rect 1156 4967 1167 4973
rect 1145 4964 1167 4967
rect 1229 4971 1243 4973
rect 1229 4965 1232 4971
rect 1239 4965 1243 4971
rect 1229 4958 1243 4965
rect 1250 4969 1269 4973
rect 1250 4961 1254 4969
rect 1263 4961 1269 4969
rect 1250 4958 1269 4961
rect 1296 4969 1307 4973
rect 1296 4962 1298 4969
rect 1306 4962 1307 4969
rect 1296 4958 1307 4962
rect 1314 4967 1336 4973
rect 1314 4961 1317 4967
rect 1325 4961 1336 4967
rect 1314 4958 1336 4961
rect 1432 4971 1446 4973
rect 1432 4965 1435 4971
rect 1442 4965 1446 4971
rect 1432 4958 1446 4965
rect 1453 4969 1472 4973
rect 1453 4961 1457 4969
rect 1466 4961 1472 4969
rect 1453 4958 1472 4961
rect 1499 4969 1510 4973
rect 1499 4962 1501 4969
rect 1509 4962 1510 4969
rect 1499 4958 1510 4962
rect 1517 4967 1539 4973
rect 1517 4961 1520 4967
rect 1528 4961 1539 4967
rect 1517 4958 1539 4961
rect 1619 4971 1633 4973
rect 1619 4965 1622 4971
rect 1629 4965 1633 4971
rect 1619 4958 1633 4965
rect 1640 4969 1659 4973
rect 1640 4961 1644 4969
rect 1653 4961 1659 4969
rect 1640 4958 1659 4961
rect 1686 4969 1697 4973
rect 1686 4962 1688 4969
rect 1696 4962 1697 4969
rect 1686 4958 1697 4962
rect 1704 4967 1726 4973
rect 1704 4961 1707 4967
rect 1715 4961 1726 4967
rect 1704 4958 1726 4961
rect 1800 4971 1814 4973
rect 1800 4965 1803 4971
rect 1810 4965 1814 4971
rect 1800 4958 1814 4965
rect 1821 4969 1840 4973
rect 1821 4961 1825 4969
rect 1834 4961 1840 4969
rect 1821 4958 1840 4961
rect 1867 4969 1878 4973
rect 1867 4962 1869 4969
rect 1877 4962 1878 4969
rect 1867 4958 1878 4962
rect 1885 4967 1907 4973
rect 1885 4961 1888 4967
rect 1896 4961 1907 4967
rect 1885 4958 1907 4961
rect 2186 4969 2200 4971
rect 2186 4963 2189 4969
rect 2196 4963 2200 4969
rect 2186 4956 2200 4963
rect 2207 4967 2226 4971
rect 2207 4959 2211 4967
rect 2220 4959 2226 4967
rect 2207 4956 2226 4959
rect 2253 4967 2264 4971
rect 2253 4960 2255 4967
rect 2263 4960 2264 4967
rect 2253 4956 2264 4960
rect 2271 4965 2293 4971
rect 2271 4959 2274 4965
rect 2282 4959 2293 4965
rect 2271 4956 2293 4959
rect 2357 4949 2359 4959
rect 2369 4949 2373 4959
rect 2357 4943 2373 4949
rect 2381 4956 2397 4959
rect 2381 4946 2383 4956
rect 2393 4946 2397 4956
rect 2381 4943 2397 4946
rect 389 4685 403 4687
rect 389 4679 392 4685
rect 399 4679 403 4685
rect 389 4672 403 4679
rect 410 4683 429 4687
rect 410 4675 414 4683
rect 423 4675 429 4683
rect 410 4672 429 4675
rect 456 4683 467 4687
rect 456 4676 458 4683
rect 466 4676 467 4683
rect 456 4672 467 4676
rect 475 4681 496 4687
rect 475 4675 477 4681
rect 485 4675 496 4681
rect 475 4672 496 4675
rect 560 4665 562 4675
rect 572 4665 576 4675
rect 560 4659 576 4665
rect 584 4672 600 4675
rect 584 4662 586 4672
rect 596 4662 600 4672
rect 584 4659 600 4662
rect 672 4681 686 4683
rect 672 4675 675 4681
rect 682 4675 686 4681
rect 672 4668 686 4675
rect 693 4679 712 4683
rect 693 4671 697 4679
rect 706 4671 712 4679
rect 693 4668 712 4671
rect 739 4679 750 4683
rect 739 4672 741 4679
rect 749 4672 750 4679
rect 739 4668 750 4672
rect 757 4677 779 4683
rect 757 4671 760 4677
rect 768 4671 779 4677
rect 935 4673 946 4675
rect 757 4668 779 4671
rect 843 4661 845 4671
rect 855 4661 859 4671
rect 843 4655 859 4661
rect 867 4668 883 4671
rect 867 4658 869 4668
rect 879 4658 883 4668
rect 935 4667 937 4673
rect 943 4667 946 4673
rect 935 4664 946 4667
rect 952 4670 968 4675
rect 952 4664 956 4670
rect 962 4664 968 4670
rect 973 4670 987 4675
rect 973 4664 977 4670
rect 983 4664 987 4670
rect 993 4670 1006 4675
rect 993 4664 997 4670
rect 1003 4664 1006 4670
rect 1025 4673 1038 4675
rect 1025 4667 1028 4673
rect 1034 4667 1038 4673
rect 1025 4664 1038 4667
rect 1044 4671 1058 4675
rect 1044 4665 1046 4671
rect 1053 4665 1058 4671
rect 1044 4664 1058 4665
rect 867 4655 883 4658
rect 469 4387 483 4389
rect 469 4381 472 4387
rect 479 4381 483 4387
rect 469 4374 483 4381
rect 490 4385 509 4389
rect 490 4377 494 4385
rect 503 4377 509 4385
rect 490 4374 509 4377
rect 536 4385 547 4389
rect 536 4378 538 4385
rect 546 4378 547 4385
rect 536 4374 547 4378
rect 554 4383 576 4389
rect 554 4377 557 4383
rect 565 4377 576 4383
rect 554 4374 576 4377
rect 672 4387 686 4389
rect 672 4381 675 4387
rect 682 4381 686 4387
rect 672 4374 686 4381
rect 693 4385 712 4389
rect 693 4377 697 4385
rect 706 4377 712 4385
rect 693 4374 712 4377
rect 739 4385 750 4389
rect 739 4378 741 4385
rect 749 4378 750 4385
rect 739 4374 750 4378
rect 757 4383 779 4389
rect 757 4377 760 4383
rect 768 4377 779 4383
rect 757 4374 779 4377
rect 859 4387 873 4389
rect 859 4381 862 4387
rect 869 4381 873 4387
rect 859 4374 873 4381
rect 880 4385 899 4389
rect 880 4377 884 4385
rect 893 4377 899 4385
rect 880 4374 899 4377
rect 926 4385 937 4389
rect 926 4378 928 4385
rect 936 4378 937 4385
rect 926 4374 937 4378
rect 944 4383 966 4389
rect 944 4377 947 4383
rect 955 4377 966 4383
rect 944 4374 966 4377
rect 1040 4387 1054 4389
rect 1040 4381 1043 4387
rect 1050 4381 1054 4387
rect 1040 4374 1054 4381
rect 1061 4385 1080 4389
rect 1061 4377 1065 4385
rect 1074 4377 1080 4385
rect 1061 4374 1080 4377
rect 1107 4385 1118 4389
rect 1107 4378 1109 4385
rect 1117 4378 1118 4385
rect 1107 4374 1118 4378
rect 1125 4383 1147 4389
rect 1125 4377 1128 4383
rect 1136 4377 1147 4383
rect 1125 4374 1147 4377
rect 1209 4381 1223 4383
rect 1209 4375 1212 4381
rect 1219 4375 1223 4381
rect 1209 4368 1223 4375
rect 1230 4379 1249 4383
rect 1230 4371 1234 4379
rect 1243 4371 1249 4379
rect 1230 4368 1249 4371
rect 1276 4379 1287 4383
rect 1276 4372 1278 4379
rect 1286 4372 1287 4379
rect 1276 4368 1287 4372
rect 1294 4377 1316 4383
rect 1294 4371 1297 4377
rect 1305 4371 1316 4377
rect 1294 4368 1316 4371
rect 1412 4381 1426 4383
rect 1412 4375 1415 4381
rect 1422 4375 1426 4381
rect 1412 4368 1426 4375
rect 1433 4379 1452 4383
rect 1433 4371 1437 4379
rect 1446 4371 1452 4379
rect 1433 4368 1452 4371
rect 1479 4379 1490 4383
rect 1479 4372 1481 4379
rect 1489 4372 1490 4379
rect 1479 4368 1490 4372
rect 1497 4377 1519 4383
rect 1497 4371 1500 4377
rect 1508 4371 1519 4377
rect 1497 4368 1519 4371
rect 1599 4381 1613 4383
rect 1599 4375 1602 4381
rect 1609 4375 1613 4381
rect 1599 4368 1613 4375
rect 1620 4379 1639 4383
rect 1620 4371 1624 4379
rect 1633 4371 1639 4379
rect 1620 4368 1639 4371
rect 1666 4379 1677 4383
rect 1666 4372 1668 4379
rect 1676 4372 1677 4379
rect 1666 4368 1677 4372
rect 1684 4377 1706 4383
rect 1684 4371 1687 4377
rect 1695 4371 1706 4377
rect 1684 4368 1706 4371
rect 1780 4381 1794 4383
rect 1780 4375 1783 4381
rect 1790 4375 1794 4381
rect 1780 4368 1794 4375
rect 1801 4379 1820 4383
rect 1801 4371 1805 4379
rect 1814 4371 1820 4379
rect 1801 4368 1820 4371
rect 1847 4379 1858 4383
rect 1847 4372 1849 4379
rect 1857 4372 1858 4379
rect 1847 4368 1858 4372
rect 1865 4377 1887 4383
rect 1865 4371 1868 4377
rect 1876 4371 1887 4377
rect 1865 4368 1887 4371
rect 2187 4379 2201 4381
rect 2187 4373 2190 4379
rect 2197 4373 2201 4379
rect 2187 4366 2201 4373
rect 2208 4377 2227 4381
rect 2208 4369 2212 4377
rect 2221 4369 2227 4377
rect 2208 4366 2227 4369
rect 2254 4377 2265 4381
rect 2254 4370 2256 4377
rect 2264 4370 2265 4377
rect 2254 4366 2265 4370
rect 2272 4375 2294 4381
rect 2272 4369 2275 4375
rect 2283 4369 2294 4375
rect 2272 4366 2294 4369
rect 2358 4359 2360 4369
rect 2370 4359 2374 4369
rect 2358 4353 2374 4359
rect 2382 4366 2398 4369
rect 2382 4356 2384 4366
rect 2394 4356 2398 4366
rect 2382 4353 2398 4356
rect 369 4095 383 4097
rect 369 4089 372 4095
rect 379 4089 383 4095
rect 369 4082 383 4089
rect 390 4093 409 4097
rect 390 4085 394 4093
rect 403 4085 409 4093
rect 390 4082 409 4085
rect 436 4093 447 4097
rect 436 4086 438 4093
rect 446 4086 447 4093
rect 436 4082 447 4086
rect 455 4091 476 4097
rect 455 4085 457 4091
rect 465 4085 476 4091
rect 455 4082 476 4085
rect 540 4075 542 4085
rect 552 4075 556 4085
rect 540 4069 556 4075
rect 564 4082 580 4085
rect 564 4072 566 4082
rect 576 4072 580 4082
rect 564 4069 580 4072
rect 652 4091 666 4093
rect 652 4085 655 4091
rect 662 4085 666 4091
rect 652 4078 666 4085
rect 673 4089 692 4093
rect 673 4081 677 4089
rect 686 4081 692 4089
rect 673 4078 692 4081
rect 719 4089 730 4093
rect 719 4082 721 4089
rect 729 4082 730 4089
rect 719 4078 730 4082
rect 737 4087 759 4093
rect 737 4081 740 4087
rect 748 4081 759 4087
rect 915 4083 926 4085
rect 737 4078 759 4081
rect 823 4071 825 4081
rect 835 4071 839 4081
rect 823 4065 839 4071
rect 847 4078 863 4081
rect 847 4068 849 4078
rect 859 4068 863 4078
rect 915 4077 917 4083
rect 923 4077 926 4083
rect 915 4074 926 4077
rect 932 4080 948 4085
rect 932 4074 936 4080
rect 942 4074 948 4080
rect 953 4080 967 4085
rect 953 4074 957 4080
rect 963 4074 967 4080
rect 973 4080 986 4085
rect 973 4074 977 4080
rect 983 4074 986 4080
rect 1005 4083 1018 4085
rect 1005 4077 1008 4083
rect 1014 4077 1018 4083
rect 1005 4074 1018 4077
rect 1024 4081 1038 4085
rect 1024 4075 1026 4081
rect 1033 4075 1038 4081
rect 1024 4074 1038 4075
rect 847 4065 863 4068
rect 497 3763 511 3765
rect 497 3757 500 3763
rect 507 3757 511 3763
rect 497 3750 511 3757
rect 518 3761 537 3765
rect 518 3753 522 3761
rect 531 3753 537 3761
rect 518 3750 537 3753
rect 564 3761 575 3765
rect 564 3754 566 3761
rect 574 3754 575 3761
rect 564 3750 575 3754
rect 582 3759 604 3765
rect 582 3753 585 3759
rect 593 3753 604 3759
rect 582 3750 604 3753
rect 700 3763 714 3765
rect 700 3757 703 3763
rect 710 3757 714 3763
rect 700 3750 714 3757
rect 721 3761 740 3765
rect 721 3753 725 3761
rect 734 3753 740 3761
rect 721 3750 740 3753
rect 767 3761 778 3765
rect 767 3754 769 3761
rect 777 3754 778 3761
rect 767 3750 778 3754
rect 785 3759 807 3765
rect 785 3753 788 3759
rect 796 3753 807 3759
rect 785 3750 807 3753
rect 887 3763 901 3765
rect 887 3757 890 3763
rect 897 3757 901 3763
rect 887 3750 901 3757
rect 908 3761 927 3765
rect 908 3753 912 3761
rect 921 3753 927 3761
rect 908 3750 927 3753
rect 954 3761 965 3765
rect 954 3754 956 3761
rect 964 3754 965 3761
rect 954 3750 965 3754
rect 972 3759 994 3765
rect 972 3753 975 3759
rect 983 3753 994 3759
rect 972 3750 994 3753
rect 1068 3763 1082 3765
rect 1068 3757 1071 3763
rect 1078 3757 1082 3763
rect 1068 3750 1082 3757
rect 1089 3761 1108 3765
rect 1089 3753 1093 3761
rect 1102 3753 1108 3761
rect 1089 3750 1108 3753
rect 1135 3761 1146 3765
rect 1135 3754 1137 3761
rect 1145 3754 1146 3761
rect 1135 3750 1146 3754
rect 1153 3759 1175 3765
rect 1153 3753 1156 3759
rect 1164 3753 1175 3759
rect 1153 3750 1175 3753
rect 1237 3757 1251 3759
rect 1237 3751 1240 3757
rect 1247 3751 1251 3757
rect 1237 3744 1251 3751
rect 1258 3755 1277 3759
rect 1258 3747 1262 3755
rect 1271 3747 1277 3755
rect 1258 3744 1277 3747
rect 1304 3755 1315 3759
rect 1304 3748 1306 3755
rect 1314 3748 1315 3755
rect 1304 3744 1315 3748
rect 1322 3753 1344 3759
rect 1322 3747 1325 3753
rect 1333 3747 1344 3753
rect 1322 3744 1344 3747
rect 1440 3757 1454 3759
rect 1440 3751 1443 3757
rect 1450 3751 1454 3757
rect 1440 3744 1454 3751
rect 1461 3755 1480 3759
rect 1461 3747 1465 3755
rect 1474 3747 1480 3755
rect 1461 3744 1480 3747
rect 1507 3755 1518 3759
rect 1507 3748 1509 3755
rect 1517 3748 1518 3755
rect 1507 3744 1518 3748
rect 1525 3753 1547 3759
rect 1525 3747 1528 3753
rect 1536 3747 1547 3753
rect 1525 3744 1547 3747
rect 1627 3757 1641 3759
rect 1627 3751 1630 3757
rect 1637 3751 1641 3757
rect 1627 3744 1641 3751
rect 1648 3755 1667 3759
rect 1648 3747 1652 3755
rect 1661 3747 1667 3755
rect 1648 3744 1667 3747
rect 1694 3755 1705 3759
rect 1694 3748 1696 3755
rect 1704 3748 1705 3755
rect 1694 3744 1705 3748
rect 1712 3753 1734 3759
rect 1712 3747 1715 3753
rect 1723 3747 1734 3753
rect 1712 3744 1734 3747
rect 1808 3757 1822 3759
rect 1808 3751 1811 3757
rect 1818 3751 1822 3757
rect 1808 3744 1822 3751
rect 1829 3755 1848 3759
rect 1829 3747 1833 3755
rect 1842 3747 1848 3755
rect 1829 3744 1848 3747
rect 1875 3755 1886 3759
rect 1875 3748 1877 3755
rect 1885 3748 1886 3755
rect 1875 3744 1886 3748
rect 1893 3753 1915 3759
rect 1893 3747 1896 3753
rect 1904 3747 1915 3753
rect 1893 3744 1915 3747
rect 2188 3755 2202 3757
rect 2188 3749 2191 3755
rect 2198 3749 2202 3755
rect 2188 3742 2202 3749
rect 2209 3753 2228 3757
rect 2209 3745 2213 3753
rect 2222 3745 2228 3753
rect 2209 3742 2228 3745
rect 2255 3753 2266 3757
rect 2255 3746 2257 3753
rect 2265 3746 2266 3753
rect 2255 3742 2266 3746
rect 2273 3751 2295 3757
rect 2273 3745 2276 3751
rect 2284 3745 2295 3751
rect 2273 3742 2295 3745
rect 2359 3735 2361 3745
rect 2371 3735 2375 3745
rect 2359 3729 2375 3735
rect 2383 3742 2399 3745
rect 2383 3732 2385 3742
rect 2395 3732 2399 3742
rect 2383 3729 2399 3732
rect 2190 3579 2204 3581
rect 2190 3573 2193 3579
rect 2200 3573 2204 3579
rect 2190 3566 2204 3573
rect 2211 3577 2230 3581
rect 2211 3569 2215 3577
rect 2224 3569 2230 3577
rect 2211 3566 2230 3569
rect 2257 3577 2268 3581
rect 2257 3570 2259 3577
rect 2267 3570 2268 3577
rect 2257 3566 2268 3570
rect 2275 3575 2297 3581
rect 2275 3569 2278 3575
rect 2286 3569 2297 3575
rect 2275 3566 2297 3569
rect 2361 3559 2363 3569
rect 2373 3559 2377 3569
rect 2361 3553 2377 3559
rect 2385 3566 2401 3569
rect 2385 3556 2387 3566
rect 2397 3556 2401 3566
rect 2385 3553 2401 3556
rect 397 3471 411 3473
rect 397 3465 400 3471
rect 407 3465 411 3471
rect 397 3458 411 3465
rect 418 3469 437 3473
rect 418 3461 422 3469
rect 431 3461 437 3469
rect 418 3458 437 3461
rect 464 3469 475 3473
rect 464 3462 466 3469
rect 474 3462 475 3469
rect 464 3458 475 3462
rect 483 3467 504 3473
rect 483 3461 485 3467
rect 493 3461 504 3467
rect 483 3458 504 3461
rect 568 3451 570 3461
rect 580 3451 584 3461
rect 568 3445 584 3451
rect 592 3458 608 3461
rect 592 3448 594 3458
rect 604 3448 608 3458
rect 592 3445 608 3448
rect 680 3467 694 3469
rect 680 3461 683 3467
rect 690 3461 694 3467
rect 680 3454 694 3461
rect 701 3465 720 3469
rect 701 3457 705 3465
rect 714 3457 720 3465
rect 701 3454 720 3457
rect 747 3465 758 3469
rect 747 3458 749 3465
rect 757 3458 758 3465
rect 747 3454 758 3458
rect 765 3463 787 3469
rect 765 3457 768 3463
rect 776 3457 787 3463
rect 943 3459 954 3461
rect 765 3454 787 3457
rect 851 3447 853 3457
rect 863 3447 867 3457
rect 851 3441 867 3447
rect 875 3454 891 3457
rect 875 3444 877 3454
rect 887 3444 891 3454
rect 943 3453 945 3459
rect 951 3453 954 3459
rect 943 3450 954 3453
rect 960 3456 976 3461
rect 960 3450 964 3456
rect 970 3450 976 3456
rect 981 3456 995 3461
rect 981 3450 985 3456
rect 991 3450 995 3456
rect 1001 3456 1014 3461
rect 1001 3450 1005 3456
rect 1011 3450 1014 3456
rect 1033 3459 1046 3461
rect 1033 3453 1036 3459
rect 1042 3453 1046 3459
rect 1033 3450 1046 3453
rect 1052 3457 1066 3461
rect 1052 3451 1054 3457
rect 1061 3451 1066 3457
rect 1052 3450 1066 3451
rect 875 3441 891 3444
rect 539 3002 553 3004
rect 539 2996 542 3002
rect 549 2996 553 3002
rect 539 2989 553 2996
rect 560 3000 579 3004
rect 560 2992 564 3000
rect 573 2992 579 3000
rect 560 2989 579 2992
rect 606 3000 617 3004
rect 606 2993 608 3000
rect 616 2993 617 3000
rect 606 2989 617 2993
rect 624 2998 646 3004
rect 624 2992 627 2998
rect 635 2992 646 2998
rect 624 2989 646 2992
rect 710 2982 712 2992
rect 722 2982 726 2992
rect 710 2976 726 2982
rect 734 2989 750 2992
rect 734 2979 736 2989
rect 746 2979 750 2989
rect 734 2976 750 2979
rect 460 2908 462 2917
rect 468 2908 470 2917
rect 479 2908 483 2917
rect 1505 2913 1516 2915
rect 1505 2907 1507 2913
rect 1513 2907 1516 2913
rect 1505 2904 1516 2907
rect 1522 2910 1538 2915
rect 1522 2904 1526 2910
rect 1532 2904 1538 2910
rect 1543 2910 1557 2915
rect 1543 2904 1547 2910
rect 1553 2904 1557 2910
rect 1563 2910 1576 2915
rect 1563 2904 1567 2910
rect 1573 2904 1576 2910
rect 1582 2910 1596 2915
rect 1582 2904 1586 2910
rect 1592 2904 1596 2910
rect 1602 2910 1615 2915
rect 1602 2904 1605 2910
rect 1611 2904 1615 2910
rect 1625 2910 1639 2915
rect 1625 2904 1629 2910
rect 1635 2904 1639 2910
rect 1645 2910 1658 2915
rect 1645 2904 1648 2910
rect 1654 2904 1658 2910
rect 1668 2913 1681 2915
rect 1668 2907 1671 2913
rect 1677 2907 1681 2913
rect 1668 2904 1681 2907
rect 1687 2911 1701 2915
rect 1687 2905 1689 2911
rect 1696 2905 1701 2911
rect 1687 2904 1701 2905
rect 539 2833 553 2835
rect 539 2827 542 2833
rect 549 2827 553 2833
rect 539 2820 553 2827
rect 560 2831 579 2835
rect 560 2823 564 2831
rect 573 2823 579 2831
rect 560 2820 579 2823
rect 606 2831 617 2835
rect 606 2824 608 2831
rect 616 2824 617 2831
rect 606 2820 617 2824
rect 624 2829 646 2835
rect 624 2823 627 2829
rect 635 2823 646 2829
rect 624 2820 646 2823
rect 669 2830 680 2834
rect 669 2823 671 2830
rect 679 2823 680 2830
rect 462 2746 464 2755
rect 470 2746 472 2755
rect 481 2746 485 2755
rect 669 2819 680 2823
rect 687 2828 709 2834
rect 687 2822 690 2828
rect 698 2822 709 2828
rect 687 2819 709 2822
rect 765 2827 767 2837
rect 777 2827 781 2837
rect 765 2821 781 2827
rect 789 2834 805 2837
rect 789 2824 791 2834
rect 801 2824 805 2834
rect 789 2821 805 2824
rect 519 2674 533 2676
rect 519 2668 522 2674
rect 529 2668 533 2674
rect 519 2661 533 2668
rect 540 2672 559 2676
rect 540 2664 544 2672
rect 553 2664 559 2672
rect 540 2661 559 2664
rect 586 2672 597 2676
rect 586 2665 588 2672
rect 596 2665 597 2672
rect 586 2661 597 2665
rect 604 2670 626 2676
rect 604 2664 607 2670
rect 615 2664 626 2670
rect 604 2661 626 2664
rect 649 2671 660 2675
rect 649 2664 651 2671
rect 659 2664 660 2671
rect 461 2591 463 2600
rect 469 2591 471 2600
rect 480 2591 484 2600
rect 649 2660 660 2664
rect 667 2669 689 2675
rect 667 2663 670 2669
rect 678 2663 689 2669
rect 667 2660 689 2663
rect 717 2669 728 2673
rect 717 2662 719 2669
rect 727 2662 728 2669
rect 717 2658 728 2662
rect 735 2667 757 2673
rect 735 2661 738 2667
rect 746 2661 757 2667
rect 735 2658 757 2661
rect 785 2666 787 2676
rect 797 2666 801 2676
rect 785 2660 801 2666
rect 809 2673 825 2676
rect 809 2663 811 2673
rect 821 2663 825 2673
rect 809 2660 825 2663
rect 528 2455 542 2457
rect 528 2449 531 2455
rect 538 2449 542 2455
rect 528 2442 542 2449
rect 549 2453 568 2457
rect 549 2445 553 2453
rect 562 2445 568 2453
rect 549 2442 568 2445
rect 595 2453 606 2457
rect 595 2446 597 2453
rect 605 2446 606 2453
rect 595 2442 606 2446
rect 613 2451 635 2457
rect 613 2445 616 2451
rect 624 2445 635 2451
rect 613 2442 635 2445
rect 658 2452 669 2456
rect 658 2445 660 2452
rect 668 2445 669 2452
rect 658 2441 669 2445
rect 676 2450 698 2456
rect 676 2444 679 2450
rect 687 2444 698 2450
rect 676 2441 698 2444
rect 726 2450 737 2454
rect 726 2443 728 2450
rect 736 2443 737 2450
rect 461 2359 463 2368
rect 469 2359 471 2368
rect 480 2359 484 2368
rect 726 2439 737 2443
rect 744 2448 766 2454
rect 744 2442 747 2448
rect 755 2442 766 2448
rect 744 2439 766 2442
rect 785 2449 796 2453
rect 785 2442 787 2449
rect 795 2442 796 2449
rect 785 2438 796 2442
rect 803 2447 825 2453
rect 803 2441 806 2447
rect 814 2441 825 2447
rect 803 2438 825 2441
rect 855 2446 857 2456
rect 867 2446 871 2456
rect 855 2440 871 2446
rect 879 2453 895 2456
rect 879 2443 881 2453
rect 891 2443 895 2453
rect 879 2440 895 2443
rect 408 2065 422 2067
rect 408 2059 411 2065
rect 418 2059 422 2065
rect 408 2052 422 2059
rect 429 2063 448 2067
rect 429 2055 433 2063
rect 442 2055 448 2063
rect 429 2052 448 2055
rect 475 2063 486 2067
rect 475 2056 477 2063
rect 485 2056 486 2063
rect 475 2052 486 2056
rect 493 2061 515 2067
rect 493 2055 496 2061
rect 504 2055 515 2061
rect 493 2052 515 2055
rect 611 2065 625 2067
rect 611 2059 614 2065
rect 621 2059 625 2065
rect 611 2052 625 2059
rect 632 2063 651 2067
rect 632 2055 636 2063
rect 645 2055 651 2063
rect 632 2052 651 2055
rect 678 2063 689 2067
rect 678 2056 680 2063
rect 688 2056 689 2063
rect 678 2052 689 2056
rect 696 2061 718 2067
rect 696 2055 699 2061
rect 707 2055 718 2061
rect 696 2052 718 2055
rect 798 2065 812 2067
rect 798 2059 801 2065
rect 808 2059 812 2065
rect 798 2052 812 2059
rect 819 2063 838 2067
rect 819 2055 823 2063
rect 832 2055 838 2063
rect 819 2052 838 2055
rect 865 2063 876 2067
rect 865 2056 867 2063
rect 875 2056 876 2063
rect 865 2052 876 2056
rect 883 2061 905 2067
rect 883 2055 886 2061
rect 894 2055 905 2061
rect 883 2052 905 2055
rect 979 2065 993 2067
rect 979 2059 982 2065
rect 989 2059 993 2065
rect 979 2052 993 2059
rect 1000 2063 1019 2067
rect 1000 2055 1004 2063
rect 1013 2055 1019 2063
rect 1000 2052 1019 2055
rect 1046 2063 1057 2067
rect 1046 2056 1048 2063
rect 1056 2056 1057 2063
rect 1046 2052 1057 2056
rect 1064 2061 1086 2067
rect 1064 2055 1067 2061
rect 1075 2055 1086 2061
rect 1064 2052 1086 2055
rect 1146 2041 1148 2050
rect 1154 2041 1156 2050
rect 1165 2041 1169 2050
rect 414 1776 428 1778
rect 414 1770 417 1776
rect 424 1770 428 1776
rect 414 1763 428 1770
rect 435 1774 454 1778
rect 435 1766 439 1774
rect 448 1766 454 1774
rect 435 1763 454 1766
rect 481 1774 492 1778
rect 481 1767 483 1774
rect 491 1767 492 1774
rect 481 1763 492 1767
rect 499 1772 521 1778
rect 499 1766 502 1772
rect 510 1766 521 1772
rect 499 1763 521 1766
rect 617 1776 631 1778
rect 617 1770 620 1776
rect 627 1770 631 1776
rect 617 1763 631 1770
rect 638 1774 657 1778
rect 638 1766 642 1774
rect 651 1766 657 1774
rect 638 1763 657 1766
rect 684 1774 695 1778
rect 684 1767 686 1774
rect 694 1767 695 1774
rect 684 1763 695 1767
rect 702 1772 724 1778
rect 702 1766 705 1772
rect 713 1766 724 1772
rect 702 1763 724 1766
rect 804 1776 818 1778
rect 804 1770 807 1776
rect 814 1770 818 1776
rect 804 1763 818 1770
rect 825 1774 844 1778
rect 825 1766 829 1774
rect 838 1766 844 1774
rect 825 1763 844 1766
rect 871 1774 882 1778
rect 871 1767 873 1774
rect 881 1767 882 1774
rect 871 1763 882 1767
rect 889 1772 911 1778
rect 889 1766 892 1772
rect 900 1766 911 1772
rect 889 1763 911 1766
rect 985 1776 999 1778
rect 985 1770 988 1776
rect 995 1770 999 1776
rect 985 1763 999 1770
rect 1006 1774 1025 1778
rect 1006 1766 1010 1774
rect 1019 1766 1025 1774
rect 1006 1763 1025 1766
rect 1052 1774 1063 1778
rect 1052 1767 1054 1774
rect 1062 1767 1063 1774
rect 1052 1763 1063 1767
rect 1070 1772 1092 1778
rect 1070 1766 1073 1772
rect 1081 1766 1092 1772
rect 1070 1763 1092 1766
rect 1148 1749 1150 1758
rect 1156 1749 1158 1758
rect 1167 1749 1171 1758
rect 434 1459 448 1461
rect 434 1453 437 1459
rect 444 1453 448 1459
rect 434 1446 448 1453
rect 455 1457 474 1461
rect 455 1449 459 1457
rect 468 1449 474 1457
rect 455 1446 474 1449
rect 501 1457 512 1461
rect 501 1450 503 1457
rect 511 1450 512 1457
rect 501 1446 512 1450
rect 519 1455 541 1461
rect 519 1449 522 1455
rect 530 1449 541 1455
rect 519 1446 541 1449
rect 637 1459 651 1461
rect 637 1453 640 1459
rect 647 1453 651 1459
rect 637 1446 651 1453
rect 658 1457 677 1461
rect 658 1449 662 1457
rect 671 1449 677 1457
rect 658 1446 677 1449
rect 704 1457 715 1461
rect 704 1450 706 1457
rect 714 1450 715 1457
rect 704 1446 715 1450
rect 722 1455 744 1461
rect 722 1449 725 1455
rect 733 1449 744 1455
rect 722 1446 744 1449
rect 824 1459 838 1461
rect 824 1453 827 1459
rect 834 1453 838 1459
rect 824 1446 838 1453
rect 845 1457 864 1461
rect 845 1449 849 1457
rect 858 1449 864 1457
rect 845 1446 864 1449
rect 891 1457 902 1461
rect 891 1450 893 1457
rect 901 1450 902 1457
rect 891 1446 902 1450
rect 909 1455 931 1461
rect 909 1449 912 1455
rect 920 1449 931 1455
rect 909 1446 931 1449
rect 1005 1459 1019 1461
rect 1005 1453 1008 1459
rect 1015 1453 1019 1459
rect 1005 1446 1019 1453
rect 1026 1457 1045 1461
rect 1026 1449 1030 1457
rect 1039 1449 1045 1457
rect 1026 1446 1045 1449
rect 1072 1457 1083 1461
rect 1072 1450 1074 1457
rect 1082 1450 1083 1457
rect 1072 1446 1083 1450
rect 1090 1455 1112 1461
rect 1090 1449 1093 1455
rect 1101 1449 1112 1455
rect 1090 1446 1112 1449
rect 1173 1432 1175 1441
rect 1181 1432 1183 1441
rect 1192 1432 1196 1441
rect 432 1168 446 1170
rect 432 1162 435 1168
rect 442 1162 446 1168
rect 432 1155 446 1162
rect 453 1166 472 1170
rect 453 1158 457 1166
rect 466 1158 472 1166
rect 453 1155 472 1158
rect 499 1166 510 1170
rect 499 1159 501 1166
rect 509 1159 510 1166
rect 499 1155 510 1159
rect 517 1164 539 1170
rect 517 1158 520 1164
rect 528 1158 539 1164
rect 517 1155 539 1158
rect 635 1168 649 1170
rect 635 1162 638 1168
rect 645 1162 649 1168
rect 635 1155 649 1162
rect 656 1166 675 1170
rect 656 1158 660 1166
rect 669 1158 675 1166
rect 656 1155 675 1158
rect 702 1166 713 1170
rect 702 1159 704 1166
rect 712 1159 713 1166
rect 702 1155 713 1159
rect 720 1164 742 1170
rect 720 1158 723 1164
rect 731 1158 742 1164
rect 720 1155 742 1158
rect 822 1168 836 1170
rect 822 1162 825 1168
rect 832 1162 836 1168
rect 822 1155 836 1162
rect 843 1166 862 1170
rect 843 1158 847 1166
rect 856 1158 862 1166
rect 843 1155 862 1158
rect 889 1166 900 1170
rect 889 1159 891 1166
rect 899 1159 900 1166
rect 889 1155 900 1159
rect 907 1164 929 1170
rect 907 1158 910 1164
rect 918 1158 929 1164
rect 907 1155 929 1158
rect 1003 1168 1017 1170
rect 1003 1162 1006 1168
rect 1013 1162 1017 1168
rect 1003 1155 1017 1162
rect 1024 1166 1043 1170
rect 1024 1158 1028 1166
rect 1037 1158 1043 1166
rect 1024 1155 1043 1158
rect 1070 1166 1081 1170
rect 1070 1159 1072 1166
rect 1080 1159 1081 1166
rect 1070 1155 1081 1159
rect 1088 1164 1110 1170
rect 1088 1158 1091 1164
rect 1099 1158 1110 1164
rect 1088 1155 1110 1158
rect 1182 1141 1184 1150
rect 1190 1141 1192 1150
rect 1201 1141 1205 1150
rect 485 736 499 738
rect 485 730 488 736
rect 495 730 499 736
rect 485 723 499 730
rect 506 734 525 738
rect 506 726 510 734
rect 519 726 525 734
rect 506 723 525 726
rect 552 734 563 738
rect 552 727 554 734
rect 562 727 563 734
rect 552 723 563 727
rect 570 732 592 738
rect 570 726 573 732
rect 581 726 592 732
rect 570 723 592 726
rect 656 716 658 726
rect 668 716 672 726
rect 656 710 672 716
rect 680 723 696 726
rect 680 713 682 723
rect 692 713 696 723
rect 680 710 696 713
rect 406 642 408 651
rect 414 642 416 651
rect 425 642 429 651
rect 485 567 499 569
rect 485 561 488 567
rect 495 561 499 567
rect 485 554 499 561
rect 506 565 525 569
rect 506 557 510 565
rect 519 557 525 565
rect 506 554 525 557
rect 552 565 563 569
rect 552 558 554 565
rect 562 558 563 565
rect 552 554 563 558
rect 570 563 592 569
rect 570 557 573 563
rect 581 557 592 563
rect 570 554 592 557
rect 615 564 626 568
rect 615 557 617 564
rect 625 557 626 564
rect 408 480 410 489
rect 416 480 418 489
rect 427 480 431 489
rect 615 553 626 557
rect 633 562 655 568
rect 633 556 636 562
rect 644 556 655 562
rect 633 553 655 556
rect 711 561 713 571
rect 723 561 727 571
rect 711 555 727 561
rect 735 568 751 571
rect 735 558 737 568
rect 747 558 751 568
rect 735 555 751 558
rect 2078 2793 2092 2795
rect 2078 2787 2081 2793
rect 2088 2787 2092 2793
rect 2078 2780 2092 2787
rect 2099 2791 2118 2795
rect 2099 2783 2103 2791
rect 2112 2783 2118 2791
rect 2099 2780 2118 2783
rect 2145 2791 2156 2795
rect 2145 2784 2147 2791
rect 2155 2784 2156 2791
rect 2145 2780 2156 2784
rect 2164 2789 2185 2795
rect 2164 2783 2166 2789
rect 2174 2783 2185 2789
rect 2164 2780 2185 2783
rect 2215 2794 2229 2796
rect 2215 2788 2218 2794
rect 2225 2788 2229 2794
rect 2215 2781 2229 2788
rect 2237 2792 2255 2796
rect 2237 2784 2240 2792
rect 2249 2784 2255 2792
rect 2237 2781 2255 2784
rect 2288 2780 2290 2789
rect 2296 2780 2298 2789
rect 2307 2780 2311 2789
rect 2078 1494 2092 1496
rect 1357 1491 1371 1493
rect 1357 1485 1360 1491
rect 1367 1485 1371 1491
rect 1357 1478 1371 1485
rect 1378 1489 1397 1493
rect 1378 1481 1382 1489
rect 1391 1481 1397 1489
rect 1378 1478 1397 1481
rect 1424 1489 1435 1493
rect 1424 1482 1426 1489
rect 1434 1482 1435 1489
rect 1424 1478 1435 1482
rect 1442 1487 1464 1493
rect 1442 1481 1445 1487
rect 1453 1481 1464 1487
rect 1442 1478 1464 1481
rect 1494 1492 1508 1494
rect 1494 1486 1497 1492
rect 1504 1486 1508 1492
rect 1494 1479 1508 1486
rect 1515 1490 1534 1494
rect 1515 1482 1519 1490
rect 1528 1482 1534 1490
rect 1515 1479 1534 1482
rect 1561 1490 1572 1494
rect 1561 1483 1563 1490
rect 1571 1483 1572 1490
rect 1561 1479 1572 1483
rect 1579 1488 1601 1494
rect 1579 1482 1582 1488
rect 1590 1482 1601 1488
rect 1579 1479 1601 1482
rect 2078 1488 2081 1494
rect 2088 1488 2092 1494
rect 2078 1481 2092 1488
rect 2099 1492 2118 1496
rect 2099 1484 2103 1492
rect 2112 1484 2118 1492
rect 2099 1481 2118 1484
rect 2145 1492 2156 1496
rect 2145 1485 2147 1492
rect 2155 1485 2156 1492
rect 2145 1481 2156 1485
rect 2163 1490 2185 1496
rect 2163 1484 2166 1490
rect 2174 1484 2185 1490
rect 2163 1481 2185 1484
rect 2215 1495 2229 1497
rect 2215 1489 2218 1495
rect 2225 1489 2229 1495
rect 2215 1482 2229 1489
rect 2237 1493 2255 1497
rect 2237 1485 2240 1493
rect 2249 1485 2255 1493
rect 2237 1482 2255 1485
rect 1635 1468 1637 1477
rect 1643 1468 1645 1477
rect 1654 1468 1658 1477
rect 2288 1481 2290 1490
rect 2296 1481 2298 1490
rect 2307 1481 2311 1490
rect 465 408 479 410
rect 465 402 468 408
rect 475 402 479 408
rect 465 395 479 402
rect 486 406 505 410
rect 486 398 490 406
rect 499 398 505 406
rect 486 395 505 398
rect 532 406 543 410
rect 532 399 534 406
rect 542 399 543 406
rect 532 395 543 399
rect 550 404 572 410
rect 550 398 553 404
rect 561 398 572 404
rect 550 395 572 398
rect 595 405 606 409
rect 595 398 597 405
rect 605 398 606 405
rect 407 325 409 334
rect 415 325 417 334
rect 426 325 430 334
rect 595 394 606 398
rect 613 403 635 409
rect 613 397 616 403
rect 624 397 635 403
rect 613 394 635 397
rect 663 403 674 407
rect 663 396 665 403
rect 673 396 674 403
rect 663 392 674 396
rect 681 401 703 407
rect 681 395 684 401
rect 692 395 703 401
rect 681 392 703 395
rect 731 400 733 410
rect 743 400 747 410
rect 731 394 747 400
rect 755 407 771 410
rect 755 397 757 407
rect 767 397 771 407
rect 755 394 771 397
rect 474 189 488 191
rect 474 183 477 189
rect 484 183 488 189
rect 474 176 488 183
rect 495 187 514 191
rect 495 179 499 187
rect 508 179 514 187
rect 495 176 514 179
rect 541 187 552 191
rect 541 180 543 187
rect 551 180 552 187
rect 541 176 552 180
rect 559 185 581 191
rect 559 179 562 185
rect 570 179 581 185
rect 559 176 581 179
rect 604 186 615 190
rect 604 179 606 186
rect 614 179 615 186
rect 604 175 615 179
rect 622 184 644 190
rect 622 178 625 184
rect 633 178 644 184
rect 622 175 644 178
rect 672 184 683 188
rect 672 177 674 184
rect 682 177 683 184
rect 407 93 409 102
rect 415 93 417 102
rect 426 93 430 102
rect 672 173 683 177
rect 690 182 712 188
rect 690 176 693 182
rect 701 176 712 182
rect 690 173 712 176
rect 731 183 742 187
rect 731 176 733 183
rect 741 176 742 183
rect 731 172 742 176
rect 749 181 771 187
rect 749 175 752 181
rect 760 175 771 181
rect 749 172 771 175
rect 801 180 803 190
rect 813 180 817 190
rect 801 174 817 180
rect 825 187 841 190
rect 825 177 827 187
rect 837 177 841 187
rect 825 174 841 177
rect 5045 1033 5056 1035
rect 5045 1027 5047 1033
rect 5053 1027 5056 1033
rect 5045 1024 5056 1027
rect 5062 1030 5078 1035
rect 5062 1024 5066 1030
rect 5072 1024 5078 1030
rect 5083 1030 5097 1035
rect 5083 1024 5087 1030
rect 5093 1024 5097 1030
rect 5103 1030 5114 1035
rect 5103 1024 5104 1030
rect 5110 1024 5114 1030
rect 5124 1030 5138 1035
rect 5124 1024 5128 1030
rect 5134 1024 5138 1030
rect 5144 1030 5157 1035
rect 5144 1024 5147 1030
rect 5153 1024 5157 1030
rect 5167 1033 5180 1035
rect 5167 1027 5170 1033
rect 5176 1027 5180 1033
rect 5167 1024 5180 1027
rect 5186 1031 5200 1035
rect 5186 1025 5188 1031
rect 5195 1025 5200 1031
rect 5186 1024 5200 1025
rect 4788 996 4799 998
rect 4788 990 4790 996
rect 4796 990 4799 996
rect 4788 987 4799 990
rect 4805 993 4821 998
rect 4805 987 4809 993
rect 4815 987 4821 993
rect 4826 993 4840 998
rect 4826 987 4830 993
rect 4836 987 4840 993
rect 4846 993 4857 998
rect 4846 987 4847 993
rect 4853 987 4857 993
rect 4867 993 4881 998
rect 4867 987 4871 993
rect 4877 987 4881 993
rect 4887 993 4900 998
rect 4887 987 4890 993
rect 4896 987 4900 993
rect 4910 996 4923 998
rect 4910 990 4913 996
rect 4919 990 4923 996
rect 4910 987 4923 990
rect 4929 994 4943 998
rect 4929 988 4931 994
rect 4938 988 4943 994
rect 4929 987 4943 988
rect 4544 841 4555 843
rect 4544 835 4546 841
rect 4552 835 4555 841
rect 4544 832 4555 835
rect 4561 838 4577 843
rect 4561 832 4565 838
rect 4571 832 4577 838
rect 4582 838 4596 843
rect 4582 832 4586 838
rect 4592 832 4596 838
rect 4602 838 4613 843
rect 4602 832 4603 838
rect 4609 832 4613 838
rect 4623 838 4637 843
rect 4623 832 4627 838
rect 4633 832 4637 838
rect 4643 838 4656 843
rect 4643 832 4646 838
rect 4652 832 4656 838
rect 4666 841 4679 843
rect 4666 835 4669 841
rect 4675 835 4679 841
rect 4666 832 4679 835
rect 4685 839 4699 843
rect 4685 833 4687 839
rect 4694 833 4699 839
rect 4685 832 4699 833
rect 2078 663 2092 665
rect 2078 657 2081 663
rect 2088 657 2092 663
rect 2078 650 2092 657
rect 2099 661 2118 665
rect 2099 653 2103 661
rect 2112 653 2118 661
rect 2099 650 2118 653
rect 2145 661 2156 665
rect 2145 654 2147 661
rect 2155 654 2156 661
rect 2145 650 2156 654
rect 2163 659 2185 665
rect 2163 653 2166 659
rect 2174 653 2185 659
rect 2163 650 2185 653
rect 2215 664 2229 666
rect 2215 658 2218 664
rect 2225 658 2229 664
rect 2215 651 2229 658
rect 2237 662 2255 666
rect 2237 654 2240 662
rect 2249 654 2255 662
rect 2237 651 2255 654
rect 1565 647 1576 649
rect 1565 641 1567 647
rect 1573 641 1576 647
rect 1565 638 1576 641
rect 1582 644 1598 649
rect 1582 638 1586 644
rect 1592 638 1598 644
rect 1603 644 1617 649
rect 1603 638 1607 644
rect 1613 638 1617 644
rect 1623 644 1636 649
rect 1623 638 1627 644
rect 1633 638 1636 644
rect 1642 644 1656 649
rect 1642 638 1646 644
rect 1652 638 1656 644
rect 1662 644 1675 649
rect 1662 638 1665 644
rect 1671 638 1675 644
rect 1685 644 1699 649
rect 1685 638 1689 644
rect 1695 638 1699 644
rect 1705 644 1718 649
rect 1705 638 1708 644
rect 1714 638 1718 644
rect 1728 647 1741 649
rect 1728 641 1731 647
rect 1737 641 1741 647
rect 1728 638 1741 641
rect 1747 645 1761 649
rect 1747 639 1749 645
rect 1756 639 1761 645
rect 1747 638 1761 639
rect 2288 650 2290 659
rect 2296 650 2298 659
rect 2307 650 2311 659
rect 691 -311 705 -309
rect 691 -317 694 -311
rect 701 -317 705 -311
rect 691 -324 705 -317
rect 712 -313 731 -309
rect 712 -321 716 -313
rect 725 -321 731 -313
rect 712 -324 731 -321
rect 758 -313 769 -309
rect 758 -320 760 -313
rect 768 -320 769 -313
rect 758 -324 769 -320
rect 776 -315 798 -309
rect 776 -321 779 -315
rect 787 -321 798 -315
rect 776 -324 798 -321
rect 862 -331 864 -321
rect 874 -331 878 -321
rect 862 -337 878 -331
rect 886 -324 902 -321
rect 886 -334 888 -324
rect 898 -334 902 -324
rect 886 -337 902 -334
rect 1279 -354 1293 -352
rect 1279 -360 1282 -354
rect 1289 -360 1293 -354
rect 1279 -367 1293 -360
rect 1300 -356 1319 -352
rect 1300 -364 1304 -356
rect 1313 -364 1319 -356
rect 1300 -367 1319 -364
rect 1346 -356 1357 -352
rect 1346 -363 1348 -356
rect 1356 -363 1357 -356
rect 1346 -367 1357 -363
rect 1364 -358 1386 -352
rect 1364 -364 1367 -358
rect 1375 -364 1386 -358
rect 1364 -367 1386 -364
rect 1416 -353 1430 -351
rect 1416 -359 1419 -353
rect 1426 -359 1430 -353
rect 1416 -366 1430 -359
rect 1438 -355 1456 -351
rect 1438 -363 1441 -355
rect 1450 -363 1456 -355
rect 1438 -366 1456 -363
rect 1489 -367 1491 -358
rect 1497 -367 1499 -358
rect 1508 -367 1512 -358
rect 693 -509 707 -507
rect 693 -515 696 -509
rect 703 -515 707 -509
rect 693 -522 707 -515
rect 714 -511 733 -507
rect 714 -519 718 -511
rect 727 -519 733 -511
rect 714 -522 733 -519
rect 760 -511 771 -507
rect 760 -518 762 -511
rect 770 -518 771 -511
rect 760 -522 771 -518
rect 778 -513 800 -507
rect 778 -519 781 -513
rect 789 -519 800 -513
rect 778 -522 800 -519
rect 864 -529 866 -519
rect 876 -529 880 -519
rect 864 -535 880 -529
rect 888 -522 904 -519
rect 888 -532 890 -522
rect 900 -532 904 -522
rect 888 -535 904 -532
rect 1279 -544 1293 -542
rect 1279 -550 1282 -544
rect 1289 -550 1293 -544
rect 1279 -557 1293 -550
rect 1300 -546 1319 -542
rect 1300 -554 1304 -546
rect 1313 -554 1319 -546
rect 1300 -557 1319 -554
rect 1346 -546 1357 -542
rect 1346 -553 1348 -546
rect 1356 -553 1357 -546
rect 1346 -557 1357 -553
rect 1364 -548 1386 -542
rect 1364 -554 1367 -548
rect 1375 -554 1386 -548
rect 1364 -557 1386 -554
rect 1416 -543 1430 -541
rect 1416 -549 1419 -543
rect 1426 -549 1430 -543
rect 1416 -556 1430 -549
rect 1438 -545 1456 -541
rect 1438 -553 1441 -545
rect 1450 -553 1456 -545
rect 1438 -556 1456 -553
rect 1489 -557 1491 -548
rect 1497 -557 1499 -548
rect 1508 -557 1512 -548
rect 693 -707 707 -705
rect 693 -713 696 -707
rect 703 -713 707 -707
rect 693 -720 707 -713
rect 714 -709 733 -705
rect 714 -717 718 -709
rect 727 -717 733 -709
rect 714 -720 733 -717
rect 760 -709 771 -705
rect 760 -716 762 -709
rect 770 -716 771 -709
rect 760 -720 771 -716
rect 778 -711 800 -705
rect 778 -717 781 -711
rect 789 -717 800 -711
rect 778 -720 800 -717
rect 864 -727 866 -717
rect 876 -727 880 -717
rect 864 -733 880 -727
rect 888 -720 904 -717
rect 888 -730 890 -720
rect 900 -730 904 -720
rect 888 -733 904 -730
rect 1279 -750 1293 -748
rect 1279 -756 1282 -750
rect 1289 -756 1293 -750
rect 1279 -763 1293 -756
rect 1300 -752 1319 -748
rect 1300 -760 1304 -752
rect 1313 -760 1319 -752
rect 1300 -763 1319 -760
rect 1346 -752 1357 -748
rect 1346 -759 1348 -752
rect 1356 -759 1357 -752
rect 1346 -763 1357 -759
rect 1364 -754 1386 -748
rect 1364 -760 1367 -754
rect 1375 -760 1386 -754
rect 1364 -763 1386 -760
rect 1416 -749 1430 -747
rect 1416 -755 1419 -749
rect 1426 -755 1430 -749
rect 1416 -762 1430 -755
rect 1438 -751 1456 -747
rect 1438 -759 1441 -751
rect 1450 -759 1456 -751
rect 1438 -762 1456 -759
rect 1489 -763 1491 -754
rect 1497 -763 1499 -754
rect 1508 -763 1512 -754
rect 5246 660 5257 662
rect 5246 654 5248 660
rect 5254 654 5257 660
rect 5246 651 5257 654
rect 5263 657 5279 662
rect 5263 651 5267 657
rect 5273 651 5279 657
rect 5284 657 5298 662
rect 5284 651 5288 657
rect 5294 651 5298 657
rect 5304 657 5317 662
rect 5304 651 5308 657
rect 5314 651 5317 657
rect 5336 660 5349 662
rect 5336 654 5339 660
rect 5345 654 5349 660
rect 5336 651 5349 654
rect 5355 658 5369 662
rect 5355 652 5357 658
rect 5364 652 5369 658
rect 5355 651 5369 652
rect 693 -902 707 -900
rect 693 -908 696 -902
rect 703 -908 707 -902
rect 693 -915 707 -908
rect 714 -904 733 -900
rect 714 -912 718 -904
rect 727 -912 733 -904
rect 714 -915 733 -912
rect 760 -904 771 -900
rect 760 -911 762 -904
rect 770 -911 771 -904
rect 760 -915 771 -911
rect 778 -906 800 -900
rect 778 -912 781 -906
rect 789 -912 800 -906
rect 778 -915 800 -912
rect 864 -922 866 -912
rect 876 -922 880 -912
rect 864 -928 880 -922
rect 888 -915 904 -912
rect 888 -925 890 -915
rect 900 -925 904 -915
rect 888 -928 904 -925
rect 1279 -940 1293 -938
rect 1279 -946 1282 -940
rect 1289 -946 1293 -940
rect 1279 -953 1293 -946
rect 1300 -942 1319 -938
rect 1300 -950 1304 -942
rect 1313 -950 1319 -942
rect 1300 -953 1319 -950
rect 1346 -942 1357 -938
rect 1346 -949 1348 -942
rect 1356 -949 1357 -942
rect 1346 -953 1357 -949
rect 1364 -944 1386 -938
rect 1364 -950 1367 -944
rect 1375 -950 1386 -944
rect 1364 -953 1386 -950
rect 1416 -939 1430 -937
rect 1416 -945 1419 -939
rect 1426 -945 1430 -939
rect 1416 -952 1430 -945
rect 1438 -941 1456 -937
rect 1438 -949 1441 -941
rect 1450 -949 1456 -941
rect 1438 -952 1456 -949
rect 1489 -953 1491 -944
rect 1497 -953 1499 -944
rect 1508 -953 1512 -944
<< ndcontact >>
rect -660 5888 -652 5895
rect -638 5885 -628 5894
rect -597 5888 -589 5896
rect -574 5887 -566 5895
rect -457 5888 -449 5895
rect -435 5885 -425 5894
rect -394 5888 -386 5896
rect -371 5887 -363 5895
rect -270 5888 -262 5895
rect -248 5885 -238 5894
rect -207 5888 -199 5896
rect -184 5887 -176 5895
rect -89 5888 -81 5895
rect -67 5885 -57 5894
rect -26 5888 -18 5896
rect -3 5887 5 5895
rect -632 5541 -624 5548
rect -610 5538 -600 5547
rect -569 5541 -561 5549
rect -546 5540 -538 5548
rect -429 5541 -421 5548
rect -407 5538 -397 5547
rect -366 5541 -358 5549
rect -343 5540 -335 5548
rect -242 5541 -234 5548
rect -220 5538 -210 5547
rect -179 5541 -171 5549
rect -156 5540 -148 5548
rect -61 5541 -53 5548
rect -39 5538 -29 5547
rect 2 5541 10 5549
rect 25 5540 33 5548
rect -632 5155 -624 5162
rect -610 5152 -600 5161
rect -569 5155 -561 5163
rect -546 5154 -538 5162
rect -429 5155 -421 5162
rect -407 5152 -397 5161
rect -366 5155 -358 5163
rect -343 5154 -335 5162
rect -242 5155 -234 5162
rect -220 5152 -210 5161
rect -179 5155 -171 5163
rect -156 5154 -148 5162
rect -61 5155 -53 5162
rect -39 5152 -29 5161
rect 2 5155 10 5163
rect 25 5154 33 5162
rect -632 4731 -624 4738
rect -610 4728 -600 4737
rect -569 4731 -561 4739
rect -546 4730 -538 4738
rect -429 4731 -421 4738
rect -407 4728 -397 4737
rect -366 4731 -358 4739
rect -343 4730 -335 4738
rect -242 4731 -234 4738
rect -220 4728 -210 4737
rect -179 4731 -171 4739
rect -156 4730 -148 4738
rect -61 4731 -53 4738
rect -39 4728 -29 4737
rect 2 4731 10 4739
rect 25 4730 33 4738
rect 434 5609 442 5616
rect 456 5606 466 5615
rect 497 5609 505 5617
rect 520 5608 528 5616
rect 637 5609 645 5616
rect 659 5606 669 5615
rect 700 5609 708 5617
rect 723 5608 731 5616
rect 824 5609 832 5616
rect 846 5606 856 5615
rect 887 5609 895 5617
rect 910 5608 918 5616
rect 1005 5609 1013 5616
rect 1027 5606 1037 5615
rect 1068 5609 1076 5617
rect 1091 5608 1099 5616
rect 1174 5603 1182 5610
rect 1196 5600 1206 5609
rect 1237 5603 1245 5611
rect 1260 5602 1268 5610
rect 1377 5603 1385 5610
rect 1399 5600 1409 5609
rect 1440 5603 1448 5611
rect 1463 5602 1471 5610
rect 1564 5603 1572 5610
rect 1586 5600 1596 5609
rect 1627 5603 1635 5611
rect 1650 5602 1658 5610
rect 1745 5603 1753 5610
rect 1767 5600 1777 5609
rect 1808 5603 1816 5611
rect 1831 5602 1839 5610
rect 3032 5644 3040 5653
rect 3050 5644 3058 5653
rect 2190 5601 2198 5608
rect 2212 5598 2222 5607
rect 2253 5601 2261 5609
rect 2276 5600 2284 5608
rect 2360 5591 2370 5601
rect 2385 5592 2395 5602
rect 3303 5567 3311 5576
rect 3321 5567 3329 5576
rect 334 5317 342 5324
rect 356 5314 366 5323
rect 397 5317 405 5325
rect 420 5316 428 5324
rect 504 5307 514 5317
rect 529 5308 539 5318
rect 617 5313 625 5320
rect 639 5310 649 5319
rect 680 5313 688 5321
rect 703 5312 711 5320
rect 880 5330 886 5335
rect 899 5330 906 5336
rect 920 5330 926 5335
rect 939 5330 946 5336
rect 971 5330 977 5335
rect 989 5330 996 5336
rect 787 5303 797 5313
rect 812 5304 822 5314
rect 491 4885 499 4892
rect 513 4882 523 4891
rect 554 4885 562 4893
rect 577 4884 585 4892
rect 694 4885 702 4892
rect 716 4882 726 4891
rect 757 4885 765 4893
rect 780 4884 788 4892
rect 881 4885 889 4892
rect 903 4882 913 4891
rect 944 4885 952 4893
rect 967 4884 975 4892
rect 1062 4885 1070 4892
rect 1084 4882 1094 4891
rect 1125 4885 1133 4893
rect 1148 4884 1156 4892
rect 1231 4879 1239 4886
rect 1253 4876 1263 4885
rect 1294 4879 1302 4887
rect 1317 4878 1325 4886
rect 1434 4879 1442 4886
rect 1456 4876 1466 4885
rect 1497 4879 1505 4887
rect 1520 4878 1528 4886
rect 1621 4879 1629 4886
rect 1643 4876 1653 4885
rect 1684 4879 1692 4887
rect 1707 4878 1715 4886
rect 1802 4879 1810 4886
rect 1824 4876 1834 4885
rect 1865 4879 1873 4887
rect 1888 4878 1896 4886
rect 2188 4877 2196 4884
rect 2210 4874 2220 4883
rect 2251 4877 2259 4885
rect 2274 4876 2282 4884
rect 391 4593 399 4600
rect 413 4590 423 4599
rect 454 4593 462 4601
rect 477 4592 485 4600
rect 561 4583 571 4593
rect 586 4584 596 4594
rect 674 4589 682 4596
rect 696 4586 706 4595
rect 737 4589 745 4597
rect 760 4588 768 4596
rect 937 4606 943 4611
rect 956 4606 963 4612
rect 977 4606 983 4611
rect 996 4606 1003 4612
rect 1028 4606 1034 4611
rect 1046 4606 1053 4612
rect 844 4579 854 4589
rect 869 4580 879 4590
rect 2358 4867 2368 4877
rect 2383 4868 2393 4878
rect 471 4295 479 4302
rect 493 4292 503 4301
rect 534 4295 542 4303
rect 557 4294 565 4302
rect 674 4295 682 4302
rect 696 4292 706 4301
rect 737 4295 745 4303
rect 760 4294 768 4302
rect 861 4295 869 4302
rect 883 4292 893 4301
rect 924 4295 932 4303
rect 947 4294 955 4302
rect 1042 4295 1050 4302
rect 1064 4292 1074 4301
rect 1105 4295 1113 4303
rect 1128 4294 1136 4302
rect 1211 4289 1219 4296
rect 1233 4286 1243 4295
rect 1274 4289 1282 4297
rect 1297 4288 1305 4296
rect 1414 4289 1422 4296
rect 1436 4286 1446 4295
rect 1477 4289 1485 4297
rect 1500 4288 1508 4296
rect 1601 4289 1609 4296
rect 1623 4286 1633 4295
rect 1664 4289 1672 4297
rect 1687 4288 1695 4296
rect 1782 4289 1790 4296
rect 1804 4286 1814 4295
rect 1845 4289 1853 4297
rect 1868 4288 1876 4296
rect 2189 4287 2197 4294
rect 2211 4284 2221 4293
rect 2252 4287 2260 4295
rect 2275 4286 2283 4294
rect 371 4003 379 4010
rect 393 4000 403 4009
rect 434 4003 442 4011
rect 457 4002 465 4010
rect 541 3993 551 4003
rect 566 3994 576 4004
rect 654 3999 662 4006
rect 676 3996 686 4005
rect 717 3999 725 4007
rect 740 3998 748 4006
rect 917 4016 923 4021
rect 936 4016 943 4022
rect 957 4016 963 4021
rect 976 4016 983 4022
rect 1008 4016 1014 4021
rect 1026 4016 1033 4022
rect 824 3989 834 3999
rect 849 3990 859 4000
rect 2359 4277 2369 4287
rect 2384 4278 2394 4288
rect 499 3671 507 3678
rect 521 3668 531 3677
rect 562 3671 570 3679
rect 585 3670 593 3678
rect 702 3671 710 3678
rect 724 3668 734 3677
rect 765 3671 773 3679
rect 788 3670 796 3678
rect 889 3671 897 3678
rect 911 3668 921 3677
rect 952 3671 960 3679
rect 975 3670 983 3678
rect 1070 3671 1078 3678
rect 1092 3668 1102 3677
rect 1133 3671 1141 3679
rect 1156 3670 1164 3678
rect 1239 3665 1247 3672
rect 1261 3662 1271 3671
rect 1302 3665 1310 3673
rect 1325 3664 1333 3672
rect 1442 3665 1450 3672
rect 1464 3662 1474 3671
rect 1505 3665 1513 3673
rect 1528 3664 1536 3672
rect 1629 3665 1637 3672
rect 1651 3662 1661 3671
rect 1692 3665 1700 3673
rect 1715 3664 1723 3672
rect 1810 3665 1818 3672
rect 1832 3662 1842 3671
rect 1873 3665 1881 3673
rect 1896 3664 1904 3672
rect 2190 3663 2198 3670
rect 2212 3660 2222 3669
rect 2253 3663 2261 3671
rect 2276 3662 2284 3670
rect 2360 3653 2370 3663
rect 2385 3654 2395 3664
rect 2192 3487 2200 3494
rect 2214 3484 2224 3493
rect 2255 3487 2263 3495
rect 2278 3486 2286 3494
rect 399 3379 407 3386
rect 421 3376 431 3385
rect 462 3379 470 3387
rect 485 3378 493 3386
rect 569 3369 579 3379
rect 594 3370 604 3380
rect 2362 3477 2372 3487
rect 2387 3478 2397 3488
rect 682 3375 690 3382
rect 704 3372 714 3381
rect 745 3375 753 3383
rect 768 3374 776 3382
rect 945 3392 951 3397
rect 964 3392 971 3398
rect 985 3392 991 3397
rect 1004 3392 1011 3398
rect 1036 3392 1042 3397
rect 1054 3392 1061 3398
rect 852 3365 862 3375
rect 877 3366 887 3376
rect 541 2910 549 2917
rect 563 2907 573 2916
rect 604 2910 612 2918
rect 627 2909 635 2917
rect 711 2900 721 2910
rect 736 2901 746 2911
rect 452 2857 460 2866
rect 470 2857 478 2866
rect 1507 2846 1513 2851
rect 1526 2846 1533 2852
rect 1547 2846 1553 2851
rect 1566 2846 1573 2852
rect 1586 2845 1592 2851
rect 1605 2846 1612 2853
rect 1629 2845 1635 2851
rect 1647 2846 1654 2852
rect 1671 2846 1677 2851
rect 1689 2846 1696 2852
rect 541 2741 549 2748
rect 563 2738 573 2747
rect 604 2741 612 2749
rect 627 2740 635 2748
rect 667 2740 675 2748
rect 690 2739 698 2747
rect 766 2745 776 2755
rect 791 2746 801 2756
rect 454 2695 462 2704
rect 472 2695 480 2704
rect 521 2582 529 2589
rect 543 2579 553 2588
rect 584 2582 592 2590
rect 607 2581 615 2589
rect 647 2581 655 2589
rect 670 2580 678 2588
rect 715 2579 723 2587
rect 738 2578 746 2586
rect 786 2584 796 2594
rect 811 2585 821 2595
rect 453 2540 461 2549
rect 471 2540 479 2549
rect 530 2363 538 2370
rect 552 2360 562 2369
rect 593 2363 601 2371
rect 616 2362 624 2370
rect 656 2362 664 2370
rect 679 2361 687 2369
rect 724 2360 732 2368
rect 747 2359 755 2367
rect 783 2359 791 2367
rect 806 2358 814 2366
rect 856 2364 866 2374
rect 881 2365 891 2375
rect 453 2308 461 2317
rect 471 2308 479 2317
rect 1138 1990 1146 1999
rect 1156 1990 1164 1999
rect 410 1973 418 1980
rect 432 1970 442 1979
rect 473 1973 481 1981
rect 496 1972 504 1980
rect 613 1973 621 1980
rect 635 1970 645 1979
rect 676 1973 684 1981
rect 699 1972 707 1980
rect 800 1973 808 1980
rect 822 1970 832 1979
rect 863 1973 871 1981
rect 886 1972 894 1980
rect 981 1973 989 1980
rect 1003 1970 1013 1979
rect 1044 1973 1052 1981
rect 1067 1972 1075 1980
rect 1140 1698 1148 1707
rect 1158 1698 1166 1707
rect 416 1684 424 1691
rect 438 1681 448 1690
rect 479 1684 487 1692
rect 502 1683 510 1691
rect 619 1684 627 1691
rect 641 1681 651 1690
rect 682 1684 690 1692
rect 705 1683 713 1691
rect 806 1684 814 1691
rect 828 1681 838 1690
rect 869 1684 877 1692
rect 892 1683 900 1691
rect 987 1684 995 1691
rect 1009 1681 1019 1690
rect 1050 1684 1058 1692
rect 1073 1683 1081 1691
rect 1165 1381 1173 1390
rect 1183 1381 1191 1390
rect 436 1367 444 1374
rect 458 1364 468 1373
rect 499 1367 507 1375
rect 522 1366 530 1374
rect 639 1367 647 1374
rect 661 1364 671 1373
rect 702 1367 710 1375
rect 725 1366 733 1374
rect 826 1367 834 1374
rect 848 1364 858 1373
rect 889 1367 897 1375
rect 912 1366 920 1374
rect 1007 1367 1015 1374
rect 1029 1364 1039 1373
rect 1070 1367 1078 1375
rect 1093 1366 1101 1374
rect 1174 1090 1182 1099
rect 1192 1090 1200 1099
rect 434 1076 442 1083
rect 456 1073 466 1082
rect 497 1076 505 1084
rect 520 1075 528 1083
rect 637 1076 645 1083
rect 659 1073 669 1082
rect 700 1076 708 1084
rect 723 1075 731 1083
rect 824 1076 832 1083
rect 846 1073 856 1082
rect 887 1076 895 1084
rect 910 1075 918 1083
rect 1005 1076 1013 1083
rect 1027 1073 1037 1082
rect 1068 1076 1076 1084
rect 1091 1075 1099 1083
rect 487 644 495 651
rect 509 641 519 650
rect 550 644 558 652
rect 573 643 581 651
rect 657 634 667 644
rect 682 635 692 645
rect 398 591 406 600
rect 416 591 424 600
rect 487 475 495 482
rect 509 472 519 481
rect 550 475 558 483
rect 573 474 581 482
rect 613 474 621 482
rect 636 473 644 481
rect 712 479 722 489
rect 737 480 747 490
rect 2280 2729 2288 2738
rect 2298 2729 2306 2738
rect 2080 2701 2088 2708
rect 2102 2698 2112 2707
rect 2143 2701 2151 2709
rect 2166 2700 2174 2708
rect 2219 2701 2227 2709
rect 2239 2699 2249 2708
rect 1627 1417 1635 1426
rect 1645 1417 1653 1426
rect 2280 1430 2288 1439
rect 2298 1430 2306 1439
rect 1359 1399 1367 1406
rect 1381 1396 1391 1405
rect 1422 1399 1430 1407
rect 1445 1398 1453 1406
rect 1498 1399 1506 1407
rect 1518 1397 1528 1406
rect 1559 1400 1567 1408
rect 1582 1399 1590 1407
rect 2080 1402 2088 1409
rect 2102 1399 2112 1408
rect 2143 1402 2151 1410
rect 2166 1401 2174 1409
rect 2219 1402 2227 1410
rect 2239 1400 2249 1409
rect 400 429 408 438
rect 418 429 426 438
rect 467 316 475 323
rect 489 313 499 322
rect 530 316 538 324
rect 553 315 561 323
rect 593 315 601 323
rect 616 314 624 322
rect 661 313 669 321
rect 684 312 692 320
rect 732 318 742 328
rect 757 319 767 329
rect 399 274 407 283
rect 417 274 425 283
rect 476 97 484 104
rect 498 94 508 103
rect 539 97 547 105
rect 562 96 570 104
rect 602 96 610 104
rect 625 95 633 103
rect 670 94 678 102
rect 693 93 701 101
rect 729 93 737 101
rect 752 92 760 100
rect 802 98 812 108
rect 827 99 837 109
rect 5047 966 5053 971
rect 5066 966 5073 972
rect 5087 966 5093 971
rect 5104 966 5111 973
rect 5128 965 5134 971
rect 5146 966 5153 972
rect 5170 966 5176 971
rect 5188 966 5195 972
rect 4790 929 4796 934
rect 4809 929 4816 935
rect 4830 929 4836 934
rect 4847 929 4854 936
rect 4871 928 4877 934
rect 4889 929 4896 935
rect 4913 929 4919 934
rect 4931 929 4938 935
rect 4546 774 4552 779
rect 4565 774 4572 780
rect 4586 774 4592 779
rect 4603 774 4610 781
rect 4627 773 4633 779
rect 4645 774 4652 780
rect 4669 774 4675 779
rect 4687 774 4694 780
rect 1567 580 1573 585
rect 1586 580 1593 586
rect 1607 580 1613 585
rect 1626 580 1633 586
rect 1646 579 1652 585
rect 1665 580 1672 587
rect 1689 579 1695 585
rect 1707 580 1714 586
rect 1731 580 1737 585
rect 1749 580 1756 586
rect 2280 599 2288 608
rect 2298 599 2306 608
rect 399 42 407 51
rect 417 42 425 51
rect 2080 571 2088 578
rect 2102 568 2112 577
rect 2143 571 2151 579
rect 2166 570 2174 578
rect 2219 571 2227 579
rect 2239 569 2249 578
rect 693 -403 701 -396
rect 715 -406 725 -397
rect 756 -403 764 -395
rect 779 -404 787 -396
rect 863 -413 873 -403
rect 888 -412 898 -402
rect 1481 -418 1489 -409
rect 1499 -418 1507 -409
rect 1281 -446 1289 -439
rect 1303 -449 1313 -440
rect 1344 -446 1352 -438
rect 1367 -447 1375 -439
rect 1420 -446 1428 -438
rect 1440 -448 1450 -439
rect 695 -601 703 -594
rect 717 -604 727 -595
rect 758 -601 766 -593
rect 781 -602 789 -594
rect 865 -611 875 -601
rect 890 -610 900 -600
rect 1481 -608 1489 -599
rect 1499 -608 1507 -599
rect 1281 -636 1289 -629
rect 1303 -639 1313 -630
rect 1344 -636 1352 -628
rect 1367 -637 1375 -629
rect 1420 -636 1428 -628
rect 1440 -638 1450 -629
rect 695 -799 703 -792
rect 717 -802 727 -793
rect 758 -799 766 -791
rect 781 -800 789 -792
rect 865 -809 875 -799
rect 890 -808 900 -798
rect 5248 593 5254 598
rect 5267 593 5274 599
rect 5288 593 5294 598
rect 5307 593 5314 599
rect 5339 593 5345 598
rect 5357 593 5364 599
rect 1481 -814 1489 -805
rect 1499 -814 1507 -805
rect 1281 -842 1289 -835
rect 1303 -845 1313 -836
rect 1344 -842 1352 -834
rect 1367 -843 1375 -835
rect 1420 -842 1428 -834
rect 1440 -844 1450 -835
rect 695 -994 703 -987
rect 717 -997 727 -988
rect 758 -994 766 -986
rect 781 -995 789 -987
rect 865 -1004 875 -994
rect 890 -1003 900 -993
rect 1481 -1004 1489 -995
rect 1499 -1004 1507 -995
rect 1281 -1032 1289 -1025
rect 1303 -1035 1313 -1026
rect 1344 -1032 1352 -1024
rect 1367 -1033 1375 -1025
rect 1420 -1032 1428 -1024
rect 1440 -1034 1450 -1025
<< pdcontact >>
rect -659 5974 -652 5980
rect -637 5970 -628 5978
rect -593 5971 -585 5978
rect -574 5970 -566 5976
rect -456 5974 -449 5980
rect -434 5970 -425 5978
rect -390 5971 -382 5978
rect -371 5970 -363 5976
rect -269 5974 -262 5980
rect -247 5970 -238 5978
rect -203 5971 -195 5978
rect -184 5970 -176 5976
rect -88 5974 -81 5980
rect -66 5970 -57 5978
rect -22 5971 -14 5978
rect -3 5970 5 5976
rect -631 5627 -624 5633
rect -609 5623 -600 5631
rect -565 5624 -557 5631
rect -546 5623 -538 5629
rect -428 5627 -421 5633
rect -406 5623 -397 5631
rect -362 5624 -354 5631
rect -343 5623 -335 5629
rect -241 5627 -234 5633
rect -219 5623 -210 5631
rect -175 5624 -167 5631
rect -156 5623 -148 5629
rect -60 5627 -53 5633
rect -38 5623 -29 5631
rect 6 5624 14 5631
rect 25 5623 33 5629
rect -631 5241 -624 5247
rect -609 5237 -600 5245
rect -565 5238 -557 5245
rect -546 5237 -538 5243
rect -428 5241 -421 5247
rect -406 5237 -397 5245
rect -362 5238 -354 5245
rect -343 5237 -335 5243
rect -241 5241 -234 5247
rect -219 5237 -210 5245
rect -175 5238 -167 5245
rect -156 5237 -148 5243
rect -60 5241 -53 5247
rect -38 5237 -29 5245
rect 6 5238 14 5245
rect 25 5237 33 5243
rect -631 4817 -624 4823
rect -609 4813 -600 4821
rect -565 4814 -557 4821
rect -546 4813 -538 4819
rect -428 4817 -421 4823
rect -406 4813 -397 4821
rect -362 4814 -354 4821
rect -343 4813 -335 4819
rect -241 4817 -234 4823
rect -219 4813 -210 4821
rect -175 4814 -167 4821
rect -156 4813 -148 4819
rect -60 4817 -53 4823
rect -38 4813 -29 4821
rect 6 4814 14 4821
rect 25 4813 33 4819
rect 435 5695 442 5701
rect 457 5691 466 5699
rect 501 5692 509 5699
rect 520 5691 528 5697
rect 638 5695 645 5701
rect 660 5691 669 5699
rect 704 5692 712 5699
rect 723 5691 731 5697
rect 825 5695 832 5701
rect 847 5691 856 5699
rect 891 5692 899 5699
rect 910 5691 918 5697
rect 1006 5695 1013 5701
rect 1028 5691 1037 5699
rect 1072 5692 1080 5699
rect 1091 5691 1099 5697
rect 1175 5689 1182 5695
rect 1197 5685 1206 5693
rect 1241 5686 1249 5693
rect 1260 5685 1268 5691
rect 1378 5689 1385 5695
rect 1400 5685 1409 5693
rect 1444 5686 1452 5693
rect 1463 5685 1471 5691
rect 1565 5689 1572 5695
rect 1587 5685 1596 5693
rect 1631 5686 1639 5693
rect 1650 5685 1658 5691
rect 1746 5689 1753 5695
rect 1768 5685 1777 5693
rect 1812 5686 1820 5693
rect 1831 5685 1839 5691
rect 2191 5687 2198 5693
rect 2213 5683 2222 5691
rect 2257 5684 2265 5691
rect 2276 5683 2284 5689
rect 2361 5673 2371 5683
rect 2385 5670 2395 5680
rect 3032 5695 3040 5704
rect 3050 5695 3059 5704
rect 3303 5618 3311 5627
rect 3321 5618 3330 5627
rect 335 5403 342 5409
rect 357 5399 366 5407
rect 401 5400 409 5407
rect 420 5399 428 5405
rect 505 5389 515 5399
rect 529 5386 539 5396
rect 618 5399 625 5405
rect 640 5395 649 5403
rect 684 5396 692 5403
rect 703 5395 711 5401
rect 788 5385 798 5395
rect 812 5382 822 5392
rect 880 5391 886 5397
rect 899 5388 905 5394
rect 920 5388 926 5394
rect 940 5388 946 5394
rect 971 5391 977 5397
rect 989 5389 996 5395
rect 492 4971 499 4977
rect 514 4967 523 4975
rect 558 4968 566 4975
rect 577 4967 585 4973
rect 695 4971 702 4977
rect 717 4967 726 4975
rect 761 4968 769 4975
rect 780 4967 788 4973
rect 882 4971 889 4977
rect 904 4967 913 4975
rect 948 4968 956 4975
rect 967 4967 975 4973
rect 1063 4971 1070 4977
rect 1085 4967 1094 4975
rect 1129 4968 1137 4975
rect 1148 4967 1156 4973
rect 1232 4965 1239 4971
rect 1254 4961 1263 4969
rect 1298 4962 1306 4969
rect 1317 4961 1325 4967
rect 1435 4965 1442 4971
rect 1457 4961 1466 4969
rect 1501 4962 1509 4969
rect 1520 4961 1528 4967
rect 1622 4965 1629 4971
rect 1644 4961 1653 4969
rect 1688 4962 1696 4969
rect 1707 4961 1715 4967
rect 1803 4965 1810 4971
rect 1825 4961 1834 4969
rect 1869 4962 1877 4969
rect 1888 4961 1896 4967
rect 2189 4963 2196 4969
rect 2211 4959 2220 4967
rect 2255 4960 2263 4967
rect 2274 4959 2282 4965
rect 2359 4949 2369 4959
rect 2383 4946 2393 4956
rect 392 4679 399 4685
rect 414 4675 423 4683
rect 458 4676 466 4683
rect 477 4675 485 4681
rect 562 4665 572 4675
rect 586 4662 596 4672
rect 675 4675 682 4681
rect 697 4671 706 4679
rect 741 4672 749 4679
rect 760 4671 768 4677
rect 845 4661 855 4671
rect 869 4658 879 4668
rect 937 4667 943 4673
rect 956 4664 962 4670
rect 977 4664 983 4670
rect 997 4664 1003 4670
rect 1028 4667 1034 4673
rect 1046 4665 1053 4671
rect 472 4381 479 4387
rect 494 4377 503 4385
rect 538 4378 546 4385
rect 557 4377 565 4383
rect 675 4381 682 4387
rect 697 4377 706 4385
rect 741 4378 749 4385
rect 760 4377 768 4383
rect 862 4381 869 4387
rect 884 4377 893 4385
rect 928 4378 936 4385
rect 947 4377 955 4383
rect 1043 4381 1050 4387
rect 1065 4377 1074 4385
rect 1109 4378 1117 4385
rect 1128 4377 1136 4383
rect 1212 4375 1219 4381
rect 1234 4371 1243 4379
rect 1278 4372 1286 4379
rect 1297 4371 1305 4377
rect 1415 4375 1422 4381
rect 1437 4371 1446 4379
rect 1481 4372 1489 4379
rect 1500 4371 1508 4377
rect 1602 4375 1609 4381
rect 1624 4371 1633 4379
rect 1668 4372 1676 4379
rect 1687 4371 1695 4377
rect 1783 4375 1790 4381
rect 1805 4371 1814 4379
rect 1849 4372 1857 4379
rect 1868 4371 1876 4377
rect 2190 4373 2197 4379
rect 2212 4369 2221 4377
rect 2256 4370 2264 4377
rect 2275 4369 2283 4375
rect 2360 4359 2370 4369
rect 2384 4356 2394 4366
rect 372 4089 379 4095
rect 394 4085 403 4093
rect 438 4086 446 4093
rect 457 4085 465 4091
rect 542 4075 552 4085
rect 566 4072 576 4082
rect 655 4085 662 4091
rect 677 4081 686 4089
rect 721 4082 729 4089
rect 740 4081 748 4087
rect 825 4071 835 4081
rect 849 4068 859 4078
rect 917 4077 923 4083
rect 936 4074 942 4080
rect 957 4074 963 4080
rect 977 4074 983 4080
rect 1008 4077 1014 4083
rect 1026 4075 1033 4081
rect 500 3757 507 3763
rect 522 3753 531 3761
rect 566 3754 574 3761
rect 585 3753 593 3759
rect 703 3757 710 3763
rect 725 3753 734 3761
rect 769 3754 777 3761
rect 788 3753 796 3759
rect 890 3757 897 3763
rect 912 3753 921 3761
rect 956 3754 964 3761
rect 975 3753 983 3759
rect 1071 3757 1078 3763
rect 1093 3753 1102 3761
rect 1137 3754 1145 3761
rect 1156 3753 1164 3759
rect 1240 3751 1247 3757
rect 1262 3747 1271 3755
rect 1306 3748 1314 3755
rect 1325 3747 1333 3753
rect 1443 3751 1450 3757
rect 1465 3747 1474 3755
rect 1509 3748 1517 3755
rect 1528 3747 1536 3753
rect 1630 3751 1637 3757
rect 1652 3747 1661 3755
rect 1696 3748 1704 3755
rect 1715 3747 1723 3753
rect 1811 3751 1818 3757
rect 1833 3747 1842 3755
rect 1877 3748 1885 3755
rect 1896 3747 1904 3753
rect 2191 3749 2198 3755
rect 2213 3745 2222 3753
rect 2257 3746 2265 3753
rect 2276 3745 2284 3751
rect 2361 3735 2371 3745
rect 2385 3732 2395 3742
rect 2193 3573 2200 3579
rect 2215 3569 2224 3577
rect 2259 3570 2267 3577
rect 2278 3569 2286 3575
rect 2363 3559 2373 3569
rect 2387 3556 2397 3566
rect 400 3465 407 3471
rect 422 3461 431 3469
rect 466 3462 474 3469
rect 485 3461 493 3467
rect 570 3451 580 3461
rect 594 3448 604 3458
rect 683 3461 690 3467
rect 705 3457 714 3465
rect 749 3458 757 3465
rect 768 3457 776 3463
rect 853 3447 863 3457
rect 877 3444 887 3454
rect 945 3453 951 3459
rect 964 3450 970 3456
rect 985 3450 991 3456
rect 1005 3450 1011 3456
rect 1036 3453 1042 3459
rect 1054 3451 1061 3457
rect 542 2996 549 3002
rect 564 2992 573 3000
rect 608 2993 616 3000
rect 627 2992 635 2998
rect 712 2982 722 2992
rect 736 2979 746 2989
rect 452 2908 460 2917
rect 470 2908 479 2917
rect 1507 2907 1513 2913
rect 1526 2904 1532 2910
rect 1547 2904 1553 2910
rect 1567 2904 1573 2910
rect 1586 2904 1592 2910
rect 1605 2904 1611 2910
rect 1629 2904 1635 2910
rect 1648 2904 1654 2910
rect 1671 2907 1677 2913
rect 1689 2905 1696 2911
rect 542 2827 549 2833
rect 564 2823 573 2831
rect 608 2824 616 2831
rect 627 2823 635 2829
rect 671 2823 679 2830
rect 454 2746 462 2755
rect 472 2746 481 2755
rect 690 2822 698 2828
rect 767 2827 777 2837
rect 791 2824 801 2834
rect 522 2668 529 2674
rect 544 2664 553 2672
rect 588 2665 596 2672
rect 607 2664 615 2670
rect 651 2664 659 2671
rect 453 2591 461 2600
rect 471 2591 480 2600
rect 670 2663 678 2669
rect 719 2662 727 2669
rect 738 2661 746 2667
rect 787 2666 797 2676
rect 811 2663 821 2673
rect 531 2449 538 2455
rect 553 2445 562 2453
rect 597 2446 605 2453
rect 616 2445 624 2451
rect 660 2445 668 2452
rect 679 2444 687 2450
rect 728 2443 736 2450
rect 453 2359 461 2368
rect 471 2359 480 2368
rect 747 2442 755 2448
rect 787 2442 795 2449
rect 806 2441 814 2447
rect 857 2446 867 2456
rect 881 2443 891 2453
rect 411 2059 418 2065
rect 433 2055 442 2063
rect 477 2056 485 2063
rect 496 2055 504 2061
rect 614 2059 621 2065
rect 636 2055 645 2063
rect 680 2056 688 2063
rect 699 2055 707 2061
rect 801 2059 808 2065
rect 823 2055 832 2063
rect 867 2056 875 2063
rect 886 2055 894 2061
rect 982 2059 989 2065
rect 1004 2055 1013 2063
rect 1048 2056 1056 2063
rect 1067 2055 1075 2061
rect 1138 2041 1146 2050
rect 1156 2041 1165 2050
rect 417 1770 424 1776
rect 439 1766 448 1774
rect 483 1767 491 1774
rect 502 1766 510 1772
rect 620 1770 627 1776
rect 642 1766 651 1774
rect 686 1767 694 1774
rect 705 1766 713 1772
rect 807 1770 814 1776
rect 829 1766 838 1774
rect 873 1767 881 1774
rect 892 1766 900 1772
rect 988 1770 995 1776
rect 1010 1766 1019 1774
rect 1054 1767 1062 1774
rect 1073 1766 1081 1772
rect 1140 1749 1148 1758
rect 1158 1749 1167 1758
rect 437 1453 444 1459
rect 459 1449 468 1457
rect 503 1450 511 1457
rect 522 1449 530 1455
rect 640 1453 647 1459
rect 662 1449 671 1457
rect 706 1450 714 1457
rect 725 1449 733 1455
rect 827 1453 834 1459
rect 849 1449 858 1457
rect 893 1450 901 1457
rect 912 1449 920 1455
rect 1008 1453 1015 1459
rect 1030 1449 1039 1457
rect 1074 1450 1082 1457
rect 1093 1449 1101 1455
rect 1165 1432 1173 1441
rect 1183 1432 1192 1441
rect 435 1162 442 1168
rect 457 1158 466 1166
rect 501 1159 509 1166
rect 520 1158 528 1164
rect 638 1162 645 1168
rect 660 1158 669 1166
rect 704 1159 712 1166
rect 723 1158 731 1164
rect 825 1162 832 1168
rect 847 1158 856 1166
rect 891 1159 899 1166
rect 910 1158 918 1164
rect 1006 1162 1013 1168
rect 1028 1158 1037 1166
rect 1072 1159 1080 1166
rect 1091 1158 1099 1164
rect 1174 1141 1182 1150
rect 1192 1141 1201 1150
rect 488 730 495 736
rect 510 726 519 734
rect 554 727 562 734
rect 573 726 581 732
rect 658 716 668 726
rect 682 713 692 723
rect 398 642 406 651
rect 416 642 425 651
rect 488 561 495 567
rect 510 557 519 565
rect 554 558 562 565
rect 573 557 581 563
rect 617 557 625 564
rect 400 480 408 489
rect 418 480 427 489
rect 636 556 644 562
rect 713 561 723 571
rect 737 558 747 568
rect 2081 2787 2088 2793
rect 2103 2783 2112 2791
rect 2147 2784 2155 2791
rect 2166 2783 2174 2789
rect 2218 2788 2225 2794
rect 2240 2784 2249 2792
rect 2280 2780 2288 2789
rect 2298 2780 2307 2789
rect 1360 1485 1367 1491
rect 1382 1481 1391 1489
rect 1426 1482 1434 1489
rect 1445 1481 1453 1487
rect 1497 1486 1504 1492
rect 1519 1482 1528 1490
rect 1563 1483 1571 1490
rect 1582 1482 1590 1488
rect 2081 1488 2088 1494
rect 2103 1484 2112 1492
rect 2147 1485 2155 1492
rect 2166 1484 2174 1490
rect 2218 1489 2225 1495
rect 2240 1485 2249 1493
rect 1627 1468 1635 1477
rect 1645 1468 1654 1477
rect 2280 1481 2288 1490
rect 2298 1481 2307 1490
rect 468 402 475 408
rect 490 398 499 406
rect 534 399 542 406
rect 553 398 561 404
rect 597 398 605 405
rect 399 325 407 334
rect 417 325 426 334
rect 616 397 624 403
rect 665 396 673 403
rect 684 395 692 401
rect 733 400 743 410
rect 757 397 767 407
rect 477 183 484 189
rect 499 179 508 187
rect 543 180 551 187
rect 562 179 570 185
rect 606 179 614 186
rect 625 178 633 184
rect 674 177 682 184
rect 399 93 407 102
rect 417 93 426 102
rect 693 176 701 182
rect 733 176 741 183
rect 752 175 760 181
rect 803 180 813 190
rect 827 177 837 187
rect 5047 1027 5053 1033
rect 5066 1024 5072 1030
rect 5087 1024 5093 1030
rect 5104 1024 5110 1030
rect 5128 1024 5134 1030
rect 5147 1024 5153 1030
rect 5170 1027 5176 1033
rect 5188 1025 5195 1031
rect 4790 990 4796 996
rect 4809 987 4815 993
rect 4830 987 4836 993
rect 4847 987 4853 993
rect 4871 987 4877 993
rect 4890 987 4896 993
rect 4913 990 4919 996
rect 4931 988 4938 994
rect 4546 835 4552 841
rect 4565 832 4571 838
rect 4586 832 4592 838
rect 4603 832 4609 838
rect 4627 832 4633 838
rect 4646 832 4652 838
rect 4669 835 4675 841
rect 4687 833 4694 839
rect 2081 657 2088 663
rect 2103 653 2112 661
rect 2147 654 2155 661
rect 2166 653 2174 659
rect 2218 658 2225 664
rect 2240 654 2249 662
rect 1567 641 1573 647
rect 1586 638 1592 644
rect 1607 638 1613 644
rect 1627 638 1633 644
rect 1646 638 1652 644
rect 1665 638 1671 644
rect 1689 638 1695 644
rect 1708 638 1714 644
rect 1731 641 1737 647
rect 1749 639 1756 645
rect 2280 650 2288 659
rect 2298 650 2307 659
rect 694 -317 701 -311
rect 716 -321 725 -313
rect 760 -320 768 -313
rect 779 -321 787 -315
rect 864 -331 874 -321
rect 888 -334 898 -324
rect 1282 -360 1289 -354
rect 1304 -364 1313 -356
rect 1348 -363 1356 -356
rect 1367 -364 1375 -358
rect 1419 -359 1426 -353
rect 1441 -363 1450 -355
rect 1481 -367 1489 -358
rect 1499 -367 1508 -358
rect 696 -515 703 -509
rect 718 -519 727 -511
rect 762 -518 770 -511
rect 781 -519 789 -513
rect 866 -529 876 -519
rect 890 -532 900 -522
rect 1282 -550 1289 -544
rect 1304 -554 1313 -546
rect 1348 -553 1356 -546
rect 1367 -554 1375 -548
rect 1419 -549 1426 -543
rect 1441 -553 1450 -545
rect 1481 -557 1489 -548
rect 1499 -557 1508 -548
rect 696 -713 703 -707
rect 718 -717 727 -709
rect 762 -716 770 -709
rect 781 -717 789 -711
rect 866 -727 876 -717
rect 890 -730 900 -720
rect 1282 -756 1289 -750
rect 1304 -760 1313 -752
rect 1348 -759 1356 -752
rect 1367 -760 1375 -754
rect 1419 -755 1426 -749
rect 1441 -759 1450 -751
rect 1481 -763 1489 -754
rect 1499 -763 1508 -754
rect 5248 654 5254 660
rect 5267 651 5273 657
rect 5288 651 5294 657
rect 5308 651 5314 657
rect 5339 654 5345 660
rect 5357 652 5364 658
rect 696 -908 703 -902
rect 718 -912 727 -904
rect 762 -911 770 -904
rect 781 -912 789 -906
rect 866 -922 876 -912
rect 890 -925 900 -915
rect 1282 -946 1289 -940
rect 1304 -950 1313 -942
rect 1348 -949 1356 -942
rect 1367 -950 1375 -944
rect 1419 -945 1426 -939
rect 1441 -949 1450 -941
rect 1481 -953 1489 -944
rect 1499 -953 1508 -944
<< polysilicon >>
rect 205 6278 206 6305
rect 148 6263 169 6267
rect 148 6240 149 6263
rect 168 6240 169 6263
rect 134 6187 135 6203
rect 69 6166 86 6169
rect 85 6145 86 6166
rect -719 6039 -237 6047
rect -719 6038 -577 6039
rect -826 6027 -800 6032
rect -947 6014 -942 6026
rect -826 6026 -817 6027
rect -927 6018 -817 6026
rect -803 6018 -800 6027
rect -718 6025 -693 6027
rect -718 6019 -692 6025
rect -927 6014 -800 6018
rect -826 6012 -800 6014
rect -702 5944 -692 6019
rect -648 5982 -641 5985
rect -584 5982 -577 6038
rect -445 5982 -438 5985
rect -381 5982 -374 5985
rect -258 5982 -251 6039
rect -194 5982 -187 5985
rect -77 5982 -70 6015
rect -13 5982 -6 5985
rect -648 5944 -641 5967
rect -702 5936 -641 5944
rect -648 5897 -641 5936
rect -584 5897 -577 5967
rect -445 5897 -438 5967
rect -381 5897 -374 5967
rect -258 5897 -251 5967
rect -194 5897 -187 5967
rect -77 5897 -70 5967
rect -13 5897 -6 5967
rect -648 5838 -641 5882
rect -584 5877 -577 5882
rect -445 5838 -438 5882
rect -381 5853 -374 5882
rect -258 5878 -251 5882
rect -194 5854 -187 5882
rect -77 5878 -70 5882
rect -648 5831 -438 5838
rect -13 5835 -6 5882
rect -691 5692 -209 5700
rect -691 5691 -549 5692
rect -828 5680 -711 5681
rect -828 5671 -827 5680
rect -813 5672 -721 5680
rect -690 5678 -665 5680
rect -690 5672 -664 5678
rect -813 5671 -711 5672
rect -828 5670 -711 5671
rect -674 5597 -664 5672
rect -620 5635 -613 5638
rect -556 5635 -549 5691
rect -417 5635 -410 5638
rect -353 5635 -346 5638
rect -230 5635 -223 5692
rect -166 5635 -159 5638
rect -49 5635 -42 5668
rect 15 5635 22 5638
rect -620 5597 -613 5620
rect -674 5589 -613 5597
rect -620 5550 -613 5589
rect -556 5550 -549 5620
rect -417 5550 -410 5620
rect -353 5550 -346 5620
rect -230 5550 -223 5620
rect -166 5550 -159 5620
rect -49 5550 -42 5620
rect 15 5550 22 5620
rect -620 5491 -613 5535
rect -556 5530 -549 5535
rect -417 5491 -410 5535
rect -353 5506 -346 5535
rect -230 5531 -223 5535
rect -166 5507 -159 5535
rect -49 5531 -42 5535
rect -620 5484 -410 5491
rect 15 5488 22 5535
rect -691 5306 -209 5314
rect -691 5305 -549 5306
rect -875 5292 -665 5294
rect -875 5284 -664 5292
rect -674 5211 -664 5284
rect -620 5249 -613 5252
rect -556 5249 -549 5305
rect -417 5249 -410 5252
rect -353 5249 -346 5252
rect -230 5249 -223 5306
rect -166 5249 -159 5252
rect -49 5249 -42 5282
rect 15 5249 22 5252
rect -620 5211 -613 5234
rect -674 5203 -613 5211
rect -620 5164 -613 5203
rect -556 5164 -549 5234
rect -417 5164 -410 5234
rect -353 5164 -346 5234
rect -230 5164 -223 5234
rect -166 5164 -159 5234
rect -49 5164 -42 5234
rect 15 5164 22 5234
rect -620 5105 -613 5149
rect -556 5144 -549 5149
rect -417 5105 -410 5149
rect -353 5120 -346 5149
rect -230 5145 -223 5149
rect -166 5121 -159 5149
rect -49 5145 -42 5149
rect -620 5098 -410 5105
rect 15 5102 22 5149
rect -691 4882 -209 4890
rect -691 4881 -549 4882
rect -690 4868 -665 4870
rect -690 4862 -664 4868
rect -674 4787 -664 4862
rect -620 4825 -613 4828
rect -556 4825 -549 4881
rect -417 4825 -410 4828
rect -353 4825 -346 4828
rect -230 4825 -223 4882
rect -166 4825 -159 4828
rect -49 4825 -42 4858
rect 15 4825 22 4828
rect -620 4787 -613 4810
rect -674 4779 -613 4787
rect -620 4740 -613 4779
rect -556 4740 -549 4810
rect -417 4740 -410 4810
rect -353 4740 -346 4810
rect -230 4740 -223 4810
rect -166 4740 -159 4810
rect -49 4740 -42 4810
rect 15 4740 22 4810
rect -620 4681 -613 4725
rect -556 4720 -549 4725
rect -417 4681 -410 4725
rect -353 4696 -346 4725
rect -230 4721 -223 4725
rect -166 4697 -159 4725
rect -49 4721 -42 4725
rect -620 4674 -410 4681
rect 15 4678 22 4725
rect 69 3797 86 6145
rect 115 4456 135 6187
rect 148 4998 169 6240
rect 187 5722 206 6278
rect 510 5767 857 5768
rect 518 5760 857 5767
rect 187 5709 332 5722
rect 446 5703 453 5706
rect 510 5703 517 5756
rect 649 5703 656 5706
rect 713 5703 720 5706
rect 836 5703 843 5760
rect 1250 5754 1265 5762
rect 900 5703 907 5706
rect 1017 5703 1024 5736
rect 1081 5703 1088 5706
rect 1186 5697 1193 5700
rect 1250 5697 1257 5754
rect 1581 5762 2037 5764
rect 1276 5755 2037 5762
rect 2266 5762 2941 5772
rect 1276 5754 1597 5755
rect 1389 5697 1396 5700
rect 1453 5697 1460 5700
rect 1576 5697 1583 5754
rect 1640 5697 1647 5700
rect 1757 5697 1764 5730
rect 1821 5697 1828 5700
rect 446 5656 453 5688
rect 446 5618 453 5645
rect 510 5618 517 5688
rect 649 5618 656 5688
rect 713 5618 720 5688
rect 836 5622 843 5688
rect 836 5618 845 5622
rect 900 5618 907 5688
rect 1017 5618 1024 5688
rect 1081 5618 1088 5688
rect 1186 5645 1193 5682
rect 1186 5612 1193 5636
rect 1250 5612 1257 5682
rect 1389 5612 1396 5682
rect 1453 5612 1460 5682
rect 1576 5612 1583 5682
rect 1640 5612 1647 5682
rect 1757 5612 1764 5682
rect 1821 5612 1828 5682
rect 446 5559 453 5603
rect 510 5598 517 5603
rect 649 5559 656 5603
rect 713 5574 720 5603
rect 446 5552 656 5559
rect 582 5496 596 5552
rect 836 5512 845 5603
rect 900 5575 907 5603
rect 1017 5599 1024 5603
rect 1081 5556 1088 5603
rect 1186 5553 1193 5597
rect 1250 5592 1257 5597
rect 1389 5553 1396 5597
rect 1453 5568 1460 5597
rect 1576 5593 1583 5597
rect 1640 5569 1647 5597
rect 1757 5593 1764 5597
rect 1186 5546 1396 5553
rect 1821 5550 1828 5597
rect 747 5502 853 5512
rect 1970 5505 1993 5755
rect 2202 5695 2209 5698
rect 2266 5695 2273 5762
rect 2375 5683 2383 5689
rect 2202 5653 2209 5680
rect 2202 5610 2209 5645
rect 2266 5610 2273 5680
rect 2931 5671 2940 5762
rect 2993 5752 3088 5759
rect 2993 5671 2999 5752
rect 3042 5704 3048 5707
rect 3042 5671 3048 5695
rect 2375 5636 2383 5667
rect 2931 5665 2999 5671
rect 3022 5665 3023 5671
rect 3028 5665 3048 5671
rect 3080 5674 3088 5752
rect 3080 5667 3088 5668
rect 2932 5664 2941 5665
rect 3042 5653 3048 5665
rect 3042 5641 3048 5644
rect 2341 5635 2383 5636
rect 2351 5626 2383 5635
rect 3313 5627 3319 5630
rect 2375 5605 2383 5626
rect 2202 5591 2209 5595
rect 2266 5550 2273 5595
rect 3313 5594 3319 5618
rect 2375 5581 2383 5589
rect 3288 5588 3319 5594
rect 3313 5576 3319 5588
rect 3313 5564 3319 5567
rect 583 5489 595 5496
rect 295 5472 457 5484
rect 593 5478 595 5489
rect 749 5486 756 5502
rect 836 5495 845 5502
rect 1152 5489 1995 5505
rect 749 5472 756 5473
rect 295 5364 307 5472
rect 1153 5452 1162 5489
rect 1970 5483 1993 5489
rect 410 5443 1162 5452
rect 346 5411 353 5414
rect 410 5411 418 5443
rect 519 5399 527 5405
rect 629 5407 636 5410
rect 693 5407 700 5433
rect 346 5364 353 5396
rect 295 5351 353 5364
rect 346 5326 353 5351
rect 410 5379 418 5396
rect 410 5326 417 5379
rect 519 5352 527 5383
rect 485 5351 527 5352
rect 495 5342 527 5351
rect 519 5321 527 5342
rect 584 5352 593 5404
rect 802 5395 810 5401
rect 889 5399 895 5403
rect 930 5399 936 5403
rect 981 5399 987 5403
rect 629 5353 636 5392
rect 600 5352 636 5353
rect 584 5344 636 5352
rect 346 5307 353 5311
rect 410 5306 417 5311
rect 519 5297 527 5305
rect 546 5276 554 5342
rect 629 5322 636 5344
rect 693 5322 700 5392
rect 802 5348 810 5379
rect 768 5347 810 5348
rect 778 5338 810 5347
rect 889 5338 895 5388
rect 930 5338 936 5388
rect 981 5366 987 5388
rect 967 5360 987 5366
rect 981 5338 987 5360
rect 2261 5375 2273 5550
rect 3250 5524 3356 5534
rect 3367 5524 3369 5534
rect 802 5317 810 5338
rect 629 5303 636 5307
rect 693 5302 700 5307
rect 802 5293 810 5301
rect 889 5277 895 5327
rect 842 5276 896 5277
rect 546 5270 896 5276
rect 547 5269 896 5270
rect 930 5252 936 5327
rect 981 5322 987 5327
rect 837 5251 936 5252
rect 849 5243 936 5251
rect 849 5242 931 5243
rect 567 5043 914 5044
rect 575 5036 914 5043
rect 143 4985 391 4998
rect 143 4983 408 4985
rect 503 4979 510 4982
rect 567 4979 574 5032
rect 706 4979 713 4982
rect 770 4979 777 4982
rect 893 4979 900 5036
rect 1307 5030 1322 5038
rect 957 4979 964 4982
rect 1074 4979 1081 5012
rect 1138 4979 1145 4982
rect 1243 4973 1250 4976
rect 1307 4973 1314 5030
rect 1638 5038 2094 5040
rect 1333 5031 2094 5038
rect 1333 5030 1654 5031
rect 1446 4973 1453 4976
rect 1510 4973 1517 4976
rect 1633 4973 1640 5030
rect 1697 4973 1704 4976
rect 1814 4973 1821 5006
rect 1878 4973 1885 4976
rect 503 4932 510 4964
rect 503 4894 510 4921
rect 567 4894 574 4964
rect 706 4894 713 4964
rect 770 4894 777 4964
rect 893 4898 900 4964
rect 893 4894 902 4898
rect 957 4894 964 4964
rect 1074 4894 1081 4964
rect 1138 4894 1145 4964
rect 1243 4921 1250 4958
rect 1243 4888 1250 4912
rect 1307 4888 1314 4958
rect 1446 4888 1453 4958
rect 1510 4888 1517 4958
rect 1633 4888 1640 4958
rect 1697 4888 1704 4958
rect 1814 4888 1821 4958
rect 1878 4888 1885 4958
rect 503 4835 510 4879
rect 567 4874 574 4879
rect 706 4835 713 4879
rect 770 4850 777 4879
rect 503 4828 713 4835
rect 639 4772 653 4828
rect 893 4788 902 4879
rect 957 4851 964 4879
rect 1074 4875 1081 4879
rect 1138 4832 1145 4879
rect 1243 4829 1250 4873
rect 1307 4868 1314 4873
rect 1446 4829 1453 4873
rect 1510 4844 1517 4873
rect 1633 4869 1640 4873
rect 1697 4845 1704 4873
rect 1814 4869 1821 4873
rect 1243 4822 1453 4829
rect 1878 4826 1885 4873
rect 804 4778 910 4788
rect 2027 4781 2050 5031
rect 2261 4983 2271 5375
rect 2200 4971 2207 4974
rect 2264 4971 2271 4983
rect 2373 4959 2381 4965
rect 2200 4929 2207 4956
rect 2200 4886 2207 4921
rect 2264 4886 2271 4956
rect 2373 4912 2381 4943
rect 2339 4911 2381 4912
rect 2349 4902 2381 4911
rect 2373 4881 2381 4902
rect 2200 4867 2207 4871
rect 640 4765 652 4772
rect 352 4748 514 4760
rect 650 4754 652 4765
rect 806 4762 813 4778
rect 893 4771 902 4778
rect 1209 4765 2052 4781
rect 806 4748 813 4749
rect 352 4640 364 4748
rect 1210 4728 1219 4765
rect 2027 4759 2050 4765
rect 467 4719 1219 4728
rect 403 4687 410 4690
rect 467 4687 475 4719
rect 576 4675 584 4681
rect 686 4683 693 4686
rect 750 4683 757 4709
rect 403 4640 410 4672
rect 352 4627 410 4640
rect 403 4602 410 4627
rect 467 4655 475 4672
rect 467 4602 474 4655
rect 576 4628 584 4659
rect 542 4627 584 4628
rect 552 4618 584 4627
rect 576 4597 584 4618
rect 641 4628 650 4680
rect 859 4671 867 4677
rect 946 4675 952 4679
rect 987 4675 993 4679
rect 1038 4675 1044 4679
rect 686 4629 693 4668
rect 657 4628 693 4629
rect 641 4620 693 4628
rect 403 4583 410 4587
rect 467 4582 474 4587
rect 576 4573 584 4581
rect 603 4552 611 4618
rect 686 4598 693 4620
rect 750 4598 757 4668
rect 859 4624 867 4655
rect 825 4623 867 4624
rect 835 4614 867 4623
rect 946 4614 952 4664
rect 987 4614 993 4664
rect 1038 4642 1044 4664
rect 1024 4636 1044 4642
rect 1038 4614 1044 4636
rect 859 4593 867 4614
rect 686 4579 693 4583
rect 750 4578 757 4583
rect 859 4569 867 4577
rect 946 4553 952 4603
rect 899 4552 953 4553
rect 603 4546 953 4552
rect 604 4545 953 4546
rect 987 4528 993 4603
rect 1038 4598 1044 4603
rect 894 4527 993 4528
rect 906 4519 993 4527
rect 906 4518 988 4519
rect 134 4437 135 4456
rect 547 4453 894 4454
rect 2264 4453 2271 4871
rect 2373 4857 2381 4865
rect 555 4446 894 4453
rect 115 4434 135 4437
rect 483 4389 490 4392
rect 547 4389 554 4442
rect 686 4389 693 4392
rect 750 4389 757 4392
rect 873 4389 880 4446
rect 1287 4440 1302 4448
rect 937 4389 944 4392
rect 1054 4389 1061 4422
rect 1118 4389 1125 4392
rect 1223 4383 1230 4386
rect 1287 4383 1294 4440
rect 1618 4448 2074 4450
rect 1313 4441 2074 4448
rect 1313 4440 1634 4441
rect 1426 4383 1433 4386
rect 1490 4383 1497 4386
rect 1613 4383 1620 4440
rect 1677 4383 1684 4386
rect 1794 4383 1801 4416
rect 1858 4383 1865 4386
rect 483 4342 490 4374
rect 483 4304 490 4331
rect 547 4304 554 4374
rect 686 4304 693 4374
rect 750 4304 757 4374
rect 873 4308 880 4374
rect 873 4304 882 4308
rect 937 4304 944 4374
rect 1054 4304 1061 4374
rect 1118 4304 1125 4374
rect 1223 4331 1230 4368
rect 1223 4298 1230 4322
rect 1287 4298 1294 4368
rect 1426 4298 1433 4368
rect 1490 4298 1497 4368
rect 1613 4298 1620 4368
rect 1677 4298 1684 4368
rect 1794 4298 1801 4368
rect 1858 4298 1865 4368
rect 483 4245 490 4289
rect 547 4284 554 4289
rect 686 4245 693 4289
rect 750 4260 757 4289
rect 483 4238 693 4245
rect 619 4182 633 4238
rect 873 4198 882 4289
rect 937 4261 944 4289
rect 1054 4285 1061 4289
rect 1118 4242 1125 4289
rect 1223 4239 1230 4283
rect 1287 4278 1294 4283
rect 1426 4239 1433 4283
rect 1490 4254 1497 4283
rect 1613 4279 1620 4283
rect 1677 4255 1684 4283
rect 1794 4279 1801 4283
rect 1223 4232 1433 4239
rect 1858 4236 1865 4283
rect 784 4188 890 4198
rect 2007 4191 2030 4441
rect 2262 4393 2272 4453
rect 2201 4381 2208 4384
rect 2265 4381 2272 4393
rect 2374 4369 2382 4375
rect 2201 4339 2208 4366
rect 2201 4296 2208 4331
rect 2265 4296 2272 4366
rect 2374 4322 2382 4353
rect 2340 4321 2382 4322
rect 2350 4312 2382 4321
rect 2374 4291 2382 4312
rect 2201 4277 2208 4281
rect 620 4175 632 4182
rect 332 4158 494 4170
rect 630 4164 632 4175
rect 786 4172 793 4188
rect 873 4181 882 4188
rect 1189 4175 2032 4191
rect 786 4158 793 4159
rect 332 4050 344 4158
rect 1190 4138 1199 4175
rect 2007 4169 2030 4175
rect 447 4129 1199 4138
rect 383 4097 390 4100
rect 447 4097 455 4129
rect 556 4085 564 4091
rect 666 4093 673 4096
rect 730 4093 737 4119
rect 383 4050 390 4082
rect 332 4037 390 4050
rect 383 4012 390 4037
rect 447 4065 455 4082
rect 447 4012 454 4065
rect 556 4038 564 4069
rect 522 4037 564 4038
rect 532 4028 564 4037
rect 556 4007 564 4028
rect 621 4038 630 4090
rect 839 4081 847 4087
rect 926 4085 932 4089
rect 967 4085 973 4089
rect 1018 4085 1024 4089
rect 666 4039 673 4078
rect 637 4038 673 4039
rect 621 4030 673 4038
rect 383 3993 390 3997
rect 447 3992 454 3997
rect 556 3983 564 3991
rect 583 3962 591 4028
rect 666 4008 673 4030
rect 730 4008 737 4078
rect 839 4034 847 4065
rect 805 4033 847 4034
rect 815 4024 847 4033
rect 926 4024 932 4074
rect 967 4024 973 4074
rect 1018 4052 1024 4074
rect 1004 4046 1024 4052
rect 1018 4024 1024 4046
rect 839 4003 847 4024
rect 666 3989 673 3993
rect 730 3988 737 3993
rect 839 3979 847 3987
rect 926 3963 932 4013
rect 879 3962 933 3963
rect 583 3956 933 3962
rect 584 3955 933 3956
rect 967 3938 973 4013
rect 1018 4008 1024 4013
rect 874 3937 973 3938
rect 886 3929 973 3937
rect 886 3928 968 3929
rect 575 3829 922 3830
rect 2265 3829 2272 4281
rect 2374 4267 2382 4275
rect 583 3822 922 3829
rect 71 3784 86 3797
rect 71 3771 74 3784
rect 85 3771 86 3784
rect 511 3765 518 3768
rect 575 3765 582 3818
rect 714 3765 721 3768
rect 778 3765 785 3768
rect 901 3765 908 3822
rect 1315 3816 1330 3824
rect 965 3765 972 3768
rect 1082 3765 1089 3798
rect 1146 3765 1153 3768
rect 1251 3759 1258 3762
rect 1315 3759 1322 3816
rect 1646 3824 2102 3826
rect 1341 3817 2102 3824
rect 1341 3816 1662 3817
rect 1454 3759 1461 3762
rect 1518 3759 1525 3762
rect 1641 3759 1648 3816
rect 1705 3759 1712 3762
rect 1822 3759 1829 3792
rect 1886 3759 1893 3762
rect 511 3718 518 3750
rect 511 3680 518 3707
rect 575 3680 582 3750
rect 714 3680 721 3750
rect 778 3680 785 3750
rect 901 3684 908 3750
rect 901 3680 910 3684
rect 965 3680 972 3750
rect 1082 3680 1089 3750
rect 1146 3680 1153 3750
rect 1251 3707 1258 3744
rect 1251 3674 1258 3698
rect 1315 3674 1322 3744
rect 1454 3674 1461 3744
rect 1518 3674 1525 3744
rect 1641 3674 1648 3744
rect 1705 3674 1712 3744
rect 1822 3674 1829 3744
rect 1886 3674 1893 3744
rect 511 3621 518 3665
rect 575 3660 582 3665
rect 714 3621 721 3665
rect 778 3636 785 3665
rect 511 3614 721 3621
rect 647 3558 661 3614
rect 901 3574 910 3665
rect 965 3637 972 3665
rect 1082 3661 1089 3665
rect 1146 3618 1153 3665
rect 1251 3615 1258 3659
rect 1315 3654 1322 3659
rect 1454 3615 1461 3659
rect 1518 3630 1525 3659
rect 1641 3655 1648 3659
rect 1705 3631 1712 3659
rect 1822 3655 1829 3659
rect 1251 3608 1461 3615
rect 1886 3612 1893 3659
rect 812 3564 918 3574
rect 2035 3567 2058 3817
rect 2263 3769 2273 3829
rect 2202 3757 2209 3760
rect 2266 3757 2273 3769
rect 2375 3745 2383 3751
rect 2202 3715 2209 3742
rect 2202 3672 2209 3707
rect 2266 3672 2273 3742
rect 2375 3698 2383 3729
rect 2341 3697 2383 3698
rect 2351 3688 2383 3697
rect 2412 3690 3226 3699
rect 2375 3667 2383 3688
rect 2202 3653 2209 3657
rect 2266 3607 2273 3657
rect 2375 3643 2383 3651
rect 2265 3593 2275 3607
rect 2204 3581 2211 3584
rect 2268 3581 2275 3593
rect 648 3551 660 3558
rect 360 3534 522 3546
rect 658 3540 660 3551
rect 814 3548 821 3564
rect 901 3557 910 3564
rect 1217 3551 2060 3567
rect 2377 3569 2385 3575
rect 814 3534 821 3535
rect 360 3426 372 3534
rect 1218 3514 1227 3551
rect 2035 3545 2058 3551
rect 475 3505 1227 3514
rect 2204 3539 2211 3566
rect 411 3473 418 3476
rect 475 3473 483 3505
rect 2204 3496 2211 3531
rect 2268 3496 2275 3566
rect 2377 3522 2385 3553
rect 2343 3521 2385 3522
rect 2353 3512 2385 3521
rect 584 3461 592 3467
rect 694 3469 701 3472
rect 758 3469 765 3495
rect 2377 3491 2385 3512
rect 2204 3477 2211 3481
rect 411 3426 418 3458
rect 360 3413 418 3426
rect 411 3388 418 3413
rect 475 3441 483 3458
rect 475 3388 482 3441
rect 584 3414 592 3445
rect 550 3413 592 3414
rect 560 3404 592 3413
rect 584 3383 592 3404
rect 649 3414 658 3466
rect 867 3457 875 3463
rect 954 3461 960 3465
rect 995 3461 1001 3465
rect 1046 3461 1052 3465
rect 694 3415 701 3454
rect 665 3414 701 3415
rect 649 3406 701 3414
rect 411 3369 418 3373
rect 475 3368 482 3373
rect 584 3359 592 3367
rect 611 3338 619 3404
rect 694 3384 701 3406
rect 758 3384 765 3454
rect 867 3410 875 3441
rect 833 3409 875 3410
rect 843 3400 875 3409
rect 954 3400 960 3450
rect 995 3400 1001 3450
rect 1046 3428 1052 3450
rect 2268 3449 2275 3481
rect 2377 3467 2385 3475
rect 1032 3422 1052 3428
rect 1046 3400 1052 3422
rect 867 3379 875 3400
rect 694 3365 701 3369
rect 758 3364 765 3369
rect 867 3355 875 3363
rect 954 3339 960 3389
rect 907 3338 961 3339
rect 611 3332 961 3338
rect 612 3331 961 3332
rect 995 3314 1001 3389
rect 1046 3384 1052 3389
rect 902 3313 1001 3314
rect 914 3305 1001 3313
rect 914 3304 996 3305
rect 2155 3167 3158 3181
rect 553 3004 560 3007
rect 617 3004 624 3007
rect 726 2992 734 2998
rect 218 2957 462 2958
rect 553 2957 560 2989
rect 218 2945 560 2957
rect 218 2944 462 2945
rect 220 2928 234 2944
rect -1298 2503 -1273 2505
rect -1421 2433 -1389 2434
rect -1421 2348 -1389 2409
rect -1363 2250 -1335 2444
rect -1298 2459 -1297 2503
rect -1248 2500 -1243 2530
rect -1221 2500 -1219 2530
rect -1298 2193 -1273 2459
rect -1274 2184 -1273 2193
rect -1298 2183 -1273 2184
rect -1248 2099 -1219 2500
rect -1171 2467 -1169 2493
rect -1220 2071 -1219 2099
rect -1189 2053 -1169 2467
rect -1152 2435 -1150 2473
rect -1138 2435 -1136 2473
rect -1152 1996 -1136 2435
rect -1110 1930 -1096 2438
rect 207 1994 215 2089
rect -122 1973 -120 1994
rect -91 1973 215 1994
rect 28 1788 196 1799
rect -135 1744 101 1745
rect -135 1728 86 1744
rect -1 1576 187 1586
rect -183 1307 95 1321
rect 220 1259 233 2928
rect 462 2917 468 2920
rect 553 2919 560 2945
rect 617 2919 624 2989
rect 726 2945 734 2976
rect 692 2944 734 2945
rect 702 2935 734 2944
rect 462 2888 468 2908
rect 726 2914 734 2935
rect 2156 2973 2163 3167
rect 3251 3084 3262 5524
rect 5321 3699 5328 3739
rect 2229 3070 3264 3084
rect 1516 2915 1522 2919
rect 1557 2915 1563 2919
rect 1596 2915 1602 2919
rect 1639 2915 1645 2919
rect 1681 2915 1687 2919
rect 553 2900 560 2904
rect 467 2881 468 2888
rect 462 2866 468 2881
rect 617 2889 624 2904
rect 726 2890 734 2898
rect 1516 2893 1522 2904
rect 462 2854 468 2857
rect 1516 2854 1522 2887
rect 1557 2854 1563 2904
rect 1596 2854 1602 2904
rect 1639 2854 1645 2904
rect 1681 2882 1687 2904
rect 1667 2876 1687 2882
rect 1681 2854 1687 2876
rect 553 2835 560 2838
rect 617 2835 624 2838
rect 781 2837 789 2843
rect 1516 2838 1522 2843
rect 680 2834 687 2837
rect 247 2788 523 2789
rect 553 2788 560 2820
rect 247 2776 560 2788
rect 248 2617 261 2776
rect 464 2755 470 2758
rect 553 2750 560 2776
rect 617 2750 624 2820
rect 464 2726 470 2746
rect 680 2749 687 2819
rect 781 2790 789 2821
rect 747 2789 789 2790
rect 757 2780 789 2789
rect 1557 2793 1563 2843
rect 781 2759 789 2780
rect 553 2731 560 2735
rect 469 2719 470 2726
rect 464 2704 470 2719
rect 617 2720 624 2735
rect 781 2735 789 2743
rect 680 2716 687 2734
rect 1235 2716 1250 2719
rect 679 2706 1250 2716
rect 464 2692 470 2695
rect 533 2676 540 2679
rect 597 2676 604 2679
rect 660 2675 667 2678
rect 801 2676 809 2682
rect 533 2633 540 2661
rect 275 2617 540 2633
rect 249 1585 259 2617
rect 275 2610 288 2617
rect 275 1847 287 2610
rect 463 2600 469 2603
rect 533 2591 540 2617
rect 597 2591 604 2661
rect 728 2673 735 2676
rect 463 2571 469 2591
rect 660 2590 667 2660
rect 533 2572 540 2576
rect 468 2564 469 2571
rect 463 2549 469 2564
rect 597 2561 604 2576
rect 728 2588 735 2658
rect 801 2629 809 2660
rect 767 2628 809 2629
rect 777 2619 809 2628
rect 801 2598 809 2619
rect 660 2557 667 2575
rect 801 2574 809 2582
rect 687 2557 697 2558
rect 659 2547 697 2557
rect 728 2555 735 2573
rect 463 2537 469 2540
rect 687 2536 697 2547
rect 727 2545 748 2555
rect 763 2545 764 2555
rect 1235 2536 1250 2706
rect 1596 2629 1602 2843
rect 1596 2613 1602 2622
rect 687 2523 1250 2536
rect 542 2457 549 2460
rect 606 2457 613 2460
rect 669 2456 676 2459
rect 504 2411 509 2413
rect 357 2398 388 2411
rect 401 2410 522 2411
rect 542 2410 549 2442
rect 401 2398 549 2410
rect 357 2132 366 2398
rect 542 2372 549 2398
rect 606 2372 613 2442
rect 737 2454 744 2457
rect 463 2368 469 2371
rect 463 2339 469 2359
rect 669 2371 676 2441
rect 796 2453 803 2494
rect 871 2456 879 2462
rect 542 2353 549 2357
rect 468 2332 469 2339
rect 463 2317 469 2332
rect 606 2342 613 2357
rect 737 2369 744 2439
rect 669 2338 676 2356
rect 796 2368 803 2438
rect 871 2409 879 2440
rect 837 2408 879 2409
rect 847 2399 879 2408
rect 871 2378 879 2399
rect 696 2338 706 2339
rect 668 2328 706 2338
rect 737 2336 744 2354
rect 871 2354 879 2362
rect 796 2347 803 2353
rect 696 2317 706 2328
rect 736 2326 757 2336
rect 772 2326 773 2336
rect 1235 2317 1250 2523
rect 1264 2557 1278 2565
rect 1264 2546 1265 2557
rect 1264 2338 1278 2546
rect 1293 2507 1307 2510
rect 463 2305 469 2308
rect 696 2304 1253 2317
rect 357 2124 833 2132
rect 357 2121 493 2124
rect 357 2120 366 2121
rect 355 2096 372 2104
rect 382 2096 383 2104
rect 355 2093 383 2096
rect 373 2017 383 2093
rect 422 2067 429 2070
rect 486 2067 493 2121
rect 625 2067 632 2070
rect 689 2067 696 2070
rect 812 2067 819 2124
rect 876 2067 883 2070
rect 993 2067 1000 2100
rect 1057 2067 1064 2070
rect 422 2017 429 2052
rect 373 2009 429 2017
rect 373 2008 383 2009
rect 422 1982 429 2009
rect 486 1982 493 2052
rect 625 1982 632 2052
rect 689 1982 696 2052
rect 812 1982 819 2052
rect 876 1982 883 2052
rect 993 1982 1000 2052
rect 1057 1982 1064 2052
rect 1148 2050 1154 2053
rect 1148 2025 1154 2041
rect 1153 2016 1154 2025
rect 1148 1999 1154 2016
rect 1148 1987 1154 1990
rect 422 1923 429 1967
rect 486 1962 493 1967
rect 625 1923 632 1967
rect 689 1938 696 1967
rect 812 1963 819 1967
rect 876 1939 883 1967
rect 993 1963 1000 1967
rect 422 1916 632 1923
rect 1057 1920 1064 1967
rect 288 1835 839 1843
rect 288 1832 499 1835
rect 371 1804 389 1815
rect 379 1728 389 1804
rect 428 1778 435 1781
rect 492 1778 499 1832
rect 631 1778 638 1781
rect 695 1778 702 1781
rect 818 1778 825 1835
rect 882 1778 889 1781
rect 999 1778 1006 1811
rect 1063 1778 1070 1781
rect 428 1728 435 1763
rect 379 1720 435 1728
rect 379 1719 389 1720
rect 428 1693 435 1720
rect 492 1693 499 1763
rect 631 1693 638 1763
rect 695 1693 702 1763
rect 818 1693 825 1763
rect 882 1693 889 1763
rect 999 1693 1006 1763
rect 1063 1693 1070 1763
rect 1150 1758 1156 1761
rect 1150 1733 1156 1749
rect 1155 1724 1156 1733
rect 1150 1707 1156 1724
rect 1150 1695 1156 1698
rect 428 1634 435 1678
rect 492 1673 499 1678
rect 631 1634 638 1678
rect 695 1649 702 1678
rect 818 1674 825 1678
rect 882 1650 889 1678
rect 999 1674 1006 1678
rect 428 1627 638 1634
rect 1063 1631 1070 1678
rect 249 1529 259 1576
rect 259 1526 390 1527
rect 259 1518 859 1526
rect 259 1515 519 1518
rect 393 1488 409 1498
rect 381 1487 409 1488
rect 399 1411 409 1487
rect 448 1461 455 1464
rect 512 1461 519 1515
rect 651 1461 658 1464
rect 715 1461 722 1464
rect 838 1461 845 1518
rect 902 1461 909 1464
rect 1019 1461 1026 1494
rect 1083 1461 1090 1464
rect 448 1411 455 1446
rect 399 1403 455 1411
rect 399 1402 409 1403
rect 448 1376 455 1403
rect 512 1376 519 1446
rect 651 1376 658 1446
rect 715 1376 722 1446
rect 838 1376 845 1446
rect 902 1376 909 1446
rect 1019 1376 1026 1446
rect 1083 1376 1090 1446
rect 1175 1441 1181 1444
rect 1175 1416 1181 1432
rect 1180 1407 1181 1416
rect 1175 1390 1181 1407
rect 1175 1378 1181 1381
rect 448 1317 455 1361
rect 512 1356 519 1361
rect 651 1317 658 1361
rect 715 1332 722 1361
rect 838 1357 845 1361
rect 902 1333 909 1361
rect 1019 1357 1026 1361
rect 448 1310 658 1317
rect 1083 1314 1090 1361
rect 218 1235 233 1259
rect 218 1227 857 1235
rect 218 1224 517 1227
rect 218 1223 233 1224
rect 218 1106 232 1223
rect -38 1097 233 1106
rect 218 1001 232 1097
rect 274 1001 275 1019
rect 274 416 285 1001
rect 329 622 343 1224
rect 379 1206 407 1207
rect 379 1196 382 1206
rect 395 1196 407 1206
rect 397 1123 407 1196
rect 446 1170 453 1173
rect 510 1170 517 1224
rect 649 1170 656 1173
rect 713 1170 720 1173
rect 836 1170 843 1227
rect 900 1170 907 1173
rect 1017 1170 1024 1203
rect 1081 1170 1088 1173
rect 397 1120 421 1123
rect 446 1120 453 1155
rect 397 1112 453 1120
rect 397 1111 421 1112
rect 406 1001 421 1111
rect 446 1085 453 1112
rect 510 1085 517 1155
rect 649 1085 656 1155
rect 713 1085 720 1155
rect 836 1085 843 1155
rect 900 1085 907 1155
rect 1017 1085 1024 1155
rect 1081 1085 1088 1155
rect 1184 1150 1190 1153
rect 1184 1125 1190 1141
rect 1189 1116 1190 1125
rect 1184 1099 1190 1116
rect 1235 1125 1250 2304
rect 1264 1416 1278 2326
rect 1277 1407 1278 1416
rect 1235 1116 1236 1125
rect 1184 1087 1190 1090
rect 446 1026 453 1070
rect 510 1065 517 1070
rect 649 1026 656 1070
rect 713 1041 720 1070
rect 836 1066 843 1070
rect 900 1042 907 1070
rect 1017 1066 1024 1070
rect 446 1019 656 1026
rect 1081 1023 1088 1070
rect 499 738 506 741
rect 563 738 570 741
rect 672 726 680 732
rect 383 692 389 693
rect 383 691 408 692
rect 499 691 506 723
rect 409 679 506 691
rect 383 678 408 679
rect 383 677 389 678
rect 408 651 414 654
rect 499 653 506 679
rect 563 653 570 723
rect 672 679 680 710
rect 638 678 680 679
rect 648 669 680 678
rect 408 622 414 642
rect 672 648 680 669
rect 499 634 506 638
rect 329 615 383 622
rect 413 615 414 622
rect 408 600 414 615
rect 563 623 570 638
rect 672 624 680 632
rect 408 588 414 591
rect 499 569 506 572
rect 563 569 570 572
rect 727 571 735 577
rect 626 568 633 571
rect 384 522 469 523
rect 499 522 506 554
rect 384 510 506 522
rect 410 489 416 492
rect 499 484 506 510
rect 563 484 570 554
rect 410 460 416 480
rect 626 483 633 553
rect 727 524 735 555
rect 693 523 735 524
rect 703 514 735 523
rect 727 493 735 514
rect 499 465 506 469
rect 415 453 416 460
rect 410 438 416 453
rect 563 454 570 469
rect 727 469 735 477
rect 626 450 633 468
rect 1235 453 1250 1116
rect 1264 1016 1278 1407
rect 1293 1510 1307 2494
rect 1639 2412 1645 2843
rect 1681 2838 1687 2843
rect 2092 2795 2099 2798
rect 2156 2795 2164 2973
rect 2229 2796 2237 3070
rect 4637 2915 4643 2917
rect 2971 2903 2972 2915
rect 2982 2903 4643 2915
rect 2290 2789 2296 2792
rect 2092 2746 2099 2780
rect 2092 2710 2099 2739
rect 2156 2710 2164 2780
rect 2229 2711 2237 2781
rect 2290 2753 2296 2780
rect 2335 2757 4603 2763
rect 2295 2746 2296 2753
rect 2290 2738 2296 2746
rect 2290 2726 2296 2729
rect 2092 2691 2099 2695
rect 1508 2025 1514 2044
rect 1293 1502 1294 1510
rect 1293 1026 1307 1502
rect 1508 1604 1514 2016
rect 2156 1702 2164 2695
rect 1371 1493 1378 1496
rect 1435 1493 1442 1496
rect 1508 1494 1515 1604
rect 1572 1494 1579 1497
rect 2092 1496 2099 1499
rect 2156 1496 2163 1702
rect 2229 1497 2237 2696
rect 2926 2592 2928 2606
rect 2937 2592 4435 2606
rect 2867 2523 2869 2537
rect 2878 2523 4477 2537
rect 2290 1490 2296 1493
rect 1371 1437 1378 1478
rect 1377 1428 1378 1437
rect 1371 1408 1378 1428
rect 1435 1408 1442 1478
rect 1508 1409 1515 1479
rect 1572 1409 1579 1479
rect 1637 1477 1643 1480
rect 1637 1448 1643 1468
rect 1642 1438 1643 1448
rect 1637 1426 1643 1438
rect 2092 1447 2099 1481
rect 1637 1414 1643 1417
rect 2092 1411 2099 1440
rect 2156 1411 2163 1481
rect 2229 1462 2237 1482
rect 2229 1412 2236 1462
rect 2290 1454 2296 1481
rect 3093 1454 3403 1458
rect 2295 1447 2296 1454
rect 2290 1439 2296 1447
rect 2290 1427 2296 1430
rect 1371 1389 1378 1393
rect 1435 1320 1442 1393
rect 1508 1390 1515 1394
rect 1572 1391 1579 1394
rect 2092 1392 2099 1396
rect 1572 1339 1580 1391
rect 1579 1328 1580 1339
rect 2156 1378 2163 1396
rect 2229 1378 2236 1397
rect 1436 1124 1442 1320
rect 1436 1092 1442 1117
rect 1235 450 1251 453
rect 625 440 1251 450
rect 1235 439 1251 440
rect 410 426 416 429
rect 274 306 286 416
rect 479 410 486 413
rect 543 410 550 413
rect 606 409 613 412
rect 747 410 755 416
rect 479 367 486 395
rect 384 351 486 367
rect 409 334 415 337
rect 479 325 486 351
rect 543 325 550 395
rect 674 407 681 410
rect 274 299 364 306
rect 274 298 378 299
rect 409 305 415 325
rect 606 324 613 394
rect 479 306 486 310
rect 414 298 415 305
rect 274 293 286 298
rect 409 283 415 298
rect 543 295 550 310
rect 674 322 681 392
rect 747 363 755 394
rect 713 362 755 363
rect 723 353 755 362
rect 747 332 755 353
rect 606 291 613 309
rect 747 308 755 316
rect 633 291 643 292
rect 605 281 643 291
rect 674 289 681 307
rect 409 271 415 274
rect 633 270 643 281
rect 673 279 694 289
rect 709 279 710 289
rect 1236 270 1251 439
rect 633 257 1251 270
rect 1263 291 1279 1016
rect 1263 280 1266 291
rect 1263 266 1279 280
rect 488 191 495 194
rect 552 191 559 194
rect 615 190 622 193
rect 450 145 455 147
rect 378 144 468 145
rect 488 144 495 176
rect 378 132 495 144
rect 488 106 495 132
rect 552 106 559 176
rect 683 188 690 191
rect 409 102 415 105
rect 409 73 415 93
rect 615 105 622 175
rect 742 187 749 228
rect 817 190 825 196
rect 488 87 495 91
rect 414 66 415 73
rect 409 51 415 66
rect 552 76 559 91
rect 683 103 690 173
rect 615 72 622 90
rect 742 102 749 172
rect 817 143 825 174
rect 783 142 825 143
rect 793 133 825 142
rect 817 112 825 133
rect 642 72 652 73
rect 614 62 652 72
rect 683 70 690 88
rect 817 88 825 96
rect 742 81 749 87
rect 642 51 652 62
rect 682 60 703 70
rect 718 60 719 70
rect 1236 51 1251 257
rect 1265 72 1279 266
rect 1293 241 1308 1026
rect 2156 871 2164 1378
rect 2092 665 2099 668
rect 2156 665 2163 871
rect 2229 666 2237 1378
rect 4555 843 4561 847
rect 4596 843 4602 2757
rect 4637 843 4643 2903
rect 4881 2587 4888 2590
rect 4799 998 4805 1002
rect 4840 998 4846 1026
rect 4881 998 4887 2587
rect 5138 2537 5145 2539
rect 5138 1066 5145 2523
rect 5056 1035 5062 1039
rect 5097 1035 5103 1057
rect 5138 1035 5144 1066
rect 5180 1035 5186 1039
rect 4923 998 4929 1002
rect 4799 937 4805 987
rect 4840 937 4846 987
rect 4881 937 4887 987
rect 4923 965 4929 987
rect 5056 974 5062 1024
rect 5097 974 5103 1024
rect 5138 974 5144 1024
rect 5180 1002 5186 1024
rect 5166 996 5186 1002
rect 5180 974 5186 996
rect 4909 959 4929 965
rect 4923 937 4929 959
rect 4679 843 4685 847
rect 4555 782 4561 832
rect 4596 782 4602 832
rect 4637 782 4643 832
rect 4679 810 4685 832
rect 4665 804 4685 810
rect 4679 782 4685 804
rect 1576 649 1582 653
rect 1617 649 1623 653
rect 1656 649 1662 653
rect 1699 649 1705 653
rect 1741 649 1747 653
rect 2290 659 2296 662
rect 1576 627 1582 638
rect 1576 588 1582 621
rect 1617 588 1623 638
rect 1656 588 1662 638
rect 1699 588 1705 638
rect 1741 616 1747 638
rect 1727 610 1747 616
rect 1741 588 1747 610
rect 2092 616 2099 650
rect 2092 580 2099 609
rect 2156 580 2163 650
rect 2229 631 2237 651
rect 2229 581 2236 631
rect 2290 623 2296 650
rect 2295 616 2296 623
rect 3073 619 3827 626
rect 2290 608 2296 616
rect 2290 596 2296 599
rect 1576 572 1582 577
rect 1617 527 1623 577
rect 1656 363 1662 577
rect 1656 347 1662 356
rect 1293 228 1294 241
rect 1293 209 1308 228
rect 409 39 415 42
rect 642 38 1254 51
rect 1236 0 1251 38
rect 1265 0 1279 60
rect 1294 0 1308 209
rect 1699 146 1705 577
rect 1741 572 1747 577
rect 2092 561 2099 565
rect 2156 -217 2163 565
rect 2229 562 2236 566
rect 1349 -225 2164 -217
rect 335 -276 776 -268
rect 335 -277 623 -276
rect 335 -432 352 -277
rect 705 -309 712 -306
rect 769 -309 776 -276
rect 878 -321 886 -315
rect 705 -394 712 -324
rect 769 -394 776 -324
rect 878 -368 886 -337
rect 1293 -352 1300 -349
rect 1357 -352 1364 -225
rect 1430 -267 3203 -255
rect 3218 -267 3219 -255
rect 1430 -351 1438 -267
rect 1491 -358 1497 -355
rect 844 -369 886 -368
rect 854 -378 886 -369
rect 878 -399 886 -378
rect 398 -439 608 -438
rect 705 -439 712 -409
rect 769 -414 776 -409
rect 1293 -401 1300 -367
rect 878 -423 886 -415
rect 1293 -437 1300 -408
rect 1357 -437 1364 -367
rect 1430 -386 1438 -366
rect 1430 -421 1437 -386
rect 1491 -394 1497 -367
rect 1496 -401 1497 -394
rect 4555 -395 4561 771
rect 4596 736 4602 771
rect 4637 766 4643 771
rect 4679 766 4685 771
rect 1491 -409 1497 -401
rect 1491 -421 1497 -418
rect 1430 -436 1438 -421
rect 398 -447 713 -439
rect 398 -457 413 -447
rect 1293 -456 1300 -452
rect -88 -472 200 -458
rect 468 -466 776 -465
rect 482 -474 778 -466
rect 707 -507 714 -504
rect 771 -507 778 -474
rect -137 -528 200 -514
rect 880 -519 888 -513
rect 707 -592 714 -522
rect 771 -592 778 -522
rect 880 -566 888 -535
rect 1293 -542 1300 -539
rect 1357 -542 1364 -452
rect 1430 -541 1438 -451
rect 1491 -548 1497 -545
rect 846 -567 888 -566
rect 856 -576 888 -567
rect 880 -597 888 -576
rect 1293 -591 1300 -557
rect 485 -637 616 -636
rect 707 -637 714 -607
rect 771 -612 778 -607
rect 880 -621 888 -613
rect 1293 -627 1300 -598
rect 1357 -627 1364 -557
rect 1430 -576 1438 -556
rect 1430 -626 1437 -576
rect 1491 -584 1497 -557
rect 1496 -591 1497 -584
rect 4799 -586 4805 926
rect 4840 891 4846 926
rect 4881 921 4887 926
rect 4923 921 4929 926
rect 1491 -599 1497 -591
rect 1491 -611 1497 -608
rect 485 -645 715 -637
rect 1293 -646 1300 -642
rect 338 -672 778 -664
rect 339 -759 353 -672
rect 707 -705 714 -702
rect 771 -705 778 -672
rect 880 -717 888 -711
rect 352 -773 353 -759
rect 707 -790 714 -720
rect 771 -790 778 -720
rect 880 -764 888 -733
rect 1293 -748 1300 -745
rect 1357 -748 1364 -642
rect 1430 -718 1437 -641
rect 1430 -747 1438 -718
rect 1491 -754 1497 -751
rect 846 -765 888 -764
rect 856 -774 888 -765
rect -209 -804 -207 -790
rect -183 -804 199 -790
rect 880 -795 888 -774
rect 529 -839 530 -825
rect 707 -835 714 -805
rect 771 -810 778 -805
rect 1293 -797 1300 -763
rect 880 -819 888 -811
rect 1293 -833 1300 -804
rect 1357 -833 1364 -763
rect 1430 -782 1438 -762
rect 1430 -817 1437 -782
rect 1491 -790 1497 -763
rect 1496 -797 1497 -790
rect 5056 -788 5062 963
rect 5097 937 5103 963
rect 5138 958 5144 963
rect 5180 958 5186 963
rect 5095 626 5104 937
rect 5298 714 5304 718
rect 5321 714 5328 3690
rect 5298 708 5328 714
rect 5257 662 5263 666
rect 5298 662 5304 708
rect 5321 707 5328 708
rect 5349 662 5355 666
rect 5095 616 5104 618
rect 5257 601 5263 651
rect 5298 601 5304 651
rect 5349 629 5355 651
rect 5335 623 5355 629
rect 5349 601 5355 623
rect 1491 -805 1497 -797
rect 1491 -817 1497 -814
rect 1430 -832 1438 -817
rect 518 -858 530 -839
rect 613 -843 715 -835
rect 1293 -852 1300 -848
rect 518 -859 629 -858
rect 518 -867 778 -859
rect 707 -900 714 -897
rect 771 -900 778 -867
rect 880 -912 888 -906
rect 707 -985 714 -915
rect 771 -985 778 -915
rect 880 -959 888 -928
rect 1293 -938 1300 -935
rect 1357 -938 1364 -848
rect 1430 -937 1438 -847
rect 1491 -944 1497 -941
rect 846 -960 888 -959
rect 856 -969 888 -960
rect 880 -990 888 -969
rect 1293 -987 1300 -953
rect 707 -1030 714 -1000
rect 771 -1005 778 -1000
rect 880 -1014 888 -1006
rect 1293 -1023 1300 -994
rect 1357 -1023 1364 -953
rect 1430 -972 1438 -952
rect 1430 -1022 1437 -972
rect 1491 -980 1497 -953
rect 5257 -974 5263 590
rect 5298 585 5304 590
rect 5349 585 5355 590
rect 1496 -987 1497 -980
rect 1491 -995 1497 -987
rect 1491 -1007 1497 -1004
rect 600 -1038 601 -1030
rect 620 -1038 715 -1030
rect 1293 -1042 1300 -1038
rect 1357 -1069 1364 -1038
rect 1430 -1041 1437 -1037
<< polycontact >>
rect 182 6278 205 6311
rect 149 6240 168 6263
rect 112 6187 134 6206
rect 69 6145 85 6166
rect -730 6037 -719 6048
rect -942 6013 -927 6027
rect -817 6018 -803 6027
rect -731 6019 -718 6027
rect -77 6015 -70 6022
rect -381 5845 -374 5853
rect -194 5846 -187 5854
rect -13 5828 -6 5835
rect -702 5690 -691 5701
rect -827 5671 -813 5680
rect -721 5672 -710 5680
rect -703 5672 -690 5680
rect -49 5668 -42 5675
rect -353 5498 -346 5506
rect -166 5499 -159 5507
rect 15 5481 22 5488
rect -702 5304 -691 5315
rect -891 5283 -875 5295
rect -49 5282 -42 5289
rect -353 5112 -346 5120
rect -166 5113 -159 5121
rect 15 5095 22 5102
rect -702 4880 -691 4891
rect -703 4862 -690 4870
rect -49 4858 -42 4865
rect -353 4688 -346 4696
rect -166 4689 -159 4697
rect 15 4671 22 4678
rect 509 5756 518 5767
rect 332 5708 351 5724
rect 1017 5736 1024 5743
rect 1265 5753 1276 5763
rect 1757 5730 1764 5737
rect 446 5645 453 5656
rect 1185 5636 1194 5645
rect 713 5566 720 5574
rect 900 5567 907 5575
rect 1081 5549 1088 5556
rect 1453 5560 1460 5568
rect 1640 5561 1647 5569
rect 1821 5543 1828 5550
rect 2202 5645 2209 5653
rect 3023 5665 3028 5671
rect 3080 5668 3088 5674
rect 2340 5625 2351 5635
rect 3278 5588 3288 5594
rect 457 5472 467 5487
rect 583 5478 593 5489
rect 749 5473 756 5486
rect 693 5433 700 5439
rect 583 5404 593 5415
rect 484 5341 495 5351
rect 546 5342 554 5354
rect 767 5337 778 5347
rect 962 5360 967 5366
rect 3356 5524 3367 5534
rect 837 5239 849 5251
rect 566 5032 575 5043
rect 391 4985 409 4998
rect 1074 5012 1081 5019
rect 1322 5029 1333 5039
rect 1814 5006 1821 5013
rect 503 4921 510 4932
rect 1242 4912 1251 4921
rect 770 4842 777 4850
rect 957 4843 964 4851
rect 1138 4825 1145 4832
rect 1510 4836 1517 4844
rect 1697 4837 1704 4845
rect 1878 4819 1885 4826
rect 2200 4921 2207 4929
rect 2338 4901 2349 4911
rect 514 4748 524 4763
rect 640 4754 650 4765
rect 806 4749 813 4762
rect 750 4709 757 4715
rect 640 4680 650 4691
rect 541 4617 552 4627
rect 603 4618 611 4630
rect 824 4613 835 4623
rect 1019 4636 1024 4642
rect 894 4515 906 4527
rect 112 4437 134 4456
rect 546 4442 555 4453
rect 1054 4422 1061 4429
rect 1302 4439 1313 4449
rect 1794 4416 1801 4423
rect 483 4331 490 4342
rect 1222 4322 1231 4331
rect 750 4252 757 4260
rect 937 4253 944 4261
rect 1118 4235 1125 4242
rect 1490 4246 1497 4254
rect 1677 4247 1684 4255
rect 1858 4229 1865 4236
rect 2201 4331 2208 4339
rect 2339 4311 2350 4321
rect 494 4158 504 4173
rect 620 4164 630 4175
rect 786 4159 793 4172
rect 730 4119 737 4125
rect 620 4090 630 4101
rect 521 4027 532 4037
rect 583 4028 591 4040
rect 804 4023 815 4033
rect 999 4046 1004 4052
rect 874 3925 886 3937
rect 574 3818 583 3829
rect 74 3768 85 3784
rect 1082 3798 1089 3805
rect 1330 3815 1341 3825
rect 1822 3792 1829 3799
rect 511 3707 518 3718
rect 1250 3698 1259 3707
rect 778 3628 785 3636
rect 965 3629 972 3637
rect 1146 3611 1153 3618
rect 1518 3622 1525 3630
rect 1705 3623 1712 3631
rect 1886 3605 1893 3612
rect 2202 3707 2209 3715
rect 2340 3687 2351 3697
rect 2405 3690 2412 3699
rect 3226 3690 3236 3699
rect 522 3534 532 3549
rect 648 3540 658 3551
rect 814 3535 821 3548
rect 2204 3531 2211 3539
rect 758 3495 765 3501
rect 2342 3511 2353 3521
rect 648 3466 658 3477
rect 549 3403 560 3413
rect 611 3404 619 3416
rect 832 3399 843 3409
rect 1027 3422 1032 3428
rect 902 3301 914 3313
rect 3158 3167 3165 3183
rect -1363 2444 -1335 2464
rect -1421 2409 -1389 2433
rect -1422 2322 -1389 2348
rect -1363 2225 -1335 2250
rect -1297 2459 -1272 2503
rect -1243 2500 -1221 2530
rect -1298 2184 -1274 2193
rect -1191 2467 -1171 2495
rect -1250 2070 -1220 2099
rect -1150 2435 -1138 2473
rect -1111 2438 -1096 2469
rect -1189 2038 -1167 2053
rect -1152 1978 -1136 1996
rect 207 2089 215 2094
rect -120 1973 -91 1994
rect -1110 1903 -1096 1930
rect 14 1788 28 1799
rect 196 1788 213 1799
rect -154 1728 -135 1745
rect 86 1728 101 1744
rect -16 1576 -1 1586
rect 187 1576 199 1586
rect -207 1307 -183 1321
rect 95 1307 110 1322
rect 691 2934 702 2944
rect 5321 3690 5328 3699
rect 462 2881 467 2888
rect 617 2877 625 2889
rect 1516 2887 1522 2893
rect 1662 2876 1667 2882
rect 746 2779 757 2789
rect 1557 2782 1564 2793
rect 464 2719 469 2726
rect 617 2708 625 2720
rect 463 2564 468 2571
rect 766 2618 777 2628
rect 597 2549 605 2561
rect 748 2544 763 2555
rect 1595 2622 1602 2629
rect 795 2494 804 2504
rect 388 2398 401 2411
rect 463 2332 468 2339
rect 606 2330 614 2342
rect 836 2398 847 2408
rect 757 2325 772 2336
rect 1265 2546 1280 2557
rect 1293 2494 1309 2507
rect 1263 2326 1280 2338
rect 372 2096 382 2104
rect 993 2100 1000 2107
rect 1148 2016 1153 2025
rect 689 1930 696 1938
rect 876 1931 883 1939
rect 1057 1913 1064 1920
rect 274 1831 288 1847
rect 361 1804 371 1815
rect 999 1811 1006 1818
rect 1150 1724 1155 1733
rect 695 1641 702 1649
rect 882 1642 889 1650
rect 1063 1624 1070 1631
rect 248 1576 259 1585
rect 249 1514 259 1529
rect 380 1488 393 1498
rect 1019 1494 1026 1501
rect 1175 1407 1180 1416
rect 715 1324 722 1332
rect 902 1325 909 1333
rect 1083 1307 1090 1314
rect -49 1097 -38 1106
rect 275 1001 285 1019
rect 382 1196 395 1206
rect 1017 1203 1024 1210
rect 1184 1116 1189 1125
rect 1263 1407 1277 1416
rect 1236 1116 1250 1125
rect 713 1033 720 1041
rect 900 1034 907 1042
rect 1081 1016 1088 1023
rect 383 679 409 691
rect 637 668 648 678
rect 383 615 392 622
rect 408 615 413 622
rect 563 611 571 623
rect 364 510 384 523
rect 692 513 703 523
rect 410 453 415 460
rect 563 442 571 454
rect 2972 2903 2982 2915
rect 2092 2739 2099 2746
rect 2317 2757 2335 2763
rect 2290 2746 2295 2753
rect 1639 2401 1645 2412
rect 1507 2016 1515 2025
rect 1294 1502 1307 1510
rect 2928 2592 2937 2606
rect 4435 2592 4462 2606
rect 2869 2523 2878 2537
rect 4477 2523 4495 2537
rect 1371 1428 1377 1437
rect 1637 1438 1642 1448
rect 2092 1440 2099 1447
rect 3088 1454 3093 1458
rect 3403 1454 3407 1458
rect 2290 1447 2295 1454
rect 1572 1328 1579 1339
rect 1435 1117 1443 1124
rect 364 351 384 367
rect 364 299 378 306
rect 409 298 414 305
rect 712 352 723 362
rect 543 283 551 295
rect 694 278 709 289
rect 1266 280 1281 291
rect 741 228 750 238
rect 364 132 378 145
rect 409 66 414 73
rect 552 64 560 76
rect 782 132 793 142
rect 703 59 718 70
rect 4881 2590 4888 2604
rect 4840 1026 4846 1032
rect 5138 2523 5145 2537
rect 5161 996 5166 1002
rect 4904 959 4909 965
rect 4660 804 4665 810
rect 1576 621 1582 627
rect 1722 610 1727 616
rect 2092 609 2099 616
rect 2290 616 2295 623
rect 3063 619 3073 626
rect 3827 619 3834 626
rect 1617 516 1624 527
rect 1655 356 1662 363
rect 1294 228 1310 241
rect 1264 60 1281 72
rect 1699 135 1705 146
rect 3203 -267 3218 -255
rect 843 -379 854 -369
rect 335 -446 354 -432
rect 1293 -408 1300 -401
rect 1491 -401 1496 -394
rect 4555 -399 4561 -395
rect -118 -472 -88 -458
rect 200 -472 217 -458
rect 397 -473 413 -457
rect 468 -475 482 -466
rect -155 -528 -137 -513
rect 200 -529 219 -514
rect 845 -577 856 -567
rect 471 -645 485 -636
rect 1293 -598 1300 -591
rect 1491 -591 1496 -584
rect 4799 -590 4805 -586
rect 338 -774 352 -759
rect 845 -775 856 -765
rect -207 -805 -183 -790
rect 199 -804 233 -790
rect 518 -839 529 -825
rect 1293 -804 1300 -797
rect 1491 -797 1496 -790
rect 5095 618 5104 626
rect 5330 623 5335 629
rect 5056 -792 5062 -788
rect 600 -843 613 -835
rect 845 -970 856 -960
rect 1293 -994 1300 -987
rect 5257 -978 5263 -974
rect 1491 -987 1496 -980
rect 601 -1039 620 -1030
<< metal1 >>
rect -1471 6283 182 6307
rect -1471 5211 -1449 6283
rect 205 6283 239 6307
rect -1424 6263 167 6264
rect -1424 6240 149 6263
rect -1421 6235 -1389 6240
rect -1384 6239 167 6240
rect -1421 5594 -1388 6235
rect -1363 6203 -1257 6204
rect -1363 6188 112 6203
rect -1476 2399 -1448 5211
rect -1421 2433 -1389 5594
rect -1363 2464 -1335 6188
rect -1278 6187 112 6188
rect 134 6187 135 6203
rect -1299 6164 -1274 6165
rect -1299 6146 69 6164
rect -1299 2503 -1274 6146
rect 85 6146 87 6164
rect -793 6077 237 6095
rect -789 6052 -775 6077
rect -856 6037 -730 6052
rect -947 6027 -928 6031
rect -947 6013 -942 6027
rect -927 6013 -925 6016
rect -947 5996 -925 6013
rect -1242 5959 -1216 5960
rect -1242 5956 -1125 5959
rect -943 5956 -925 5996
rect -856 5982 -842 6037
rect -814 6027 -734 6029
rect -803 6019 -731 6027
rect -328 6022 -69 6024
rect -803 6018 -734 6019
rect -814 6016 -734 6018
rect -684 6011 -343 6021
rect -328 6015 -77 6022
rect -70 6015 -69 6022
rect -328 6014 -69 6015
rect -593 6000 -585 6011
rect -390 6000 -382 6011
rect -659 5994 -585 6000
rect -761 5982 -748 5985
rect -856 5968 -748 5982
rect -659 5980 -652 5994
rect -593 5978 -585 5994
rect -1242 5939 -925 5956
rect -1242 5938 -1125 5939
rect -943 5938 -925 5939
rect -1242 2530 -1216 5938
rect -761 5710 -748 5968
rect -456 5994 -382 6000
rect -456 5980 -449 5994
rect -637 5939 -628 5970
rect -390 5978 -382 5994
rect -574 5949 -566 5970
rect -575 5939 -566 5949
rect -637 5936 -566 5939
rect -434 5939 -425 5970
rect -371 5939 -363 5970
rect -434 5938 -363 5939
rect -327 5938 -318 6014
rect -203 6000 -195 6009
rect -22 6000 -14 6009
rect -269 5994 -195 6000
rect -269 5980 -262 5994
rect -203 5978 -195 5994
rect -637 5931 -540 5936
rect -434 5931 -318 5938
rect -88 5994 -14 6000
rect -88 5980 -81 5994
rect -247 5939 -238 5970
rect -22 5978 -14 5994
rect -184 5939 -176 5970
rect -247 5938 -176 5939
rect -66 5939 -57 5970
rect -3 5939 5 5970
rect -66 5938 5 5939
rect 17 5938 125 5940
rect -247 5931 -130 5938
rect -66 5931 125 5938
rect -574 5927 -540 5931
rect -638 5903 -589 5911
rect -660 5866 -652 5888
rect -638 5894 -628 5903
rect -597 5896 -589 5903
rect -574 5895 -566 5927
rect -551 5854 -540 5927
rect -371 5929 -318 5931
rect -184 5929 -130 5931
rect -435 5903 -386 5911
rect -457 5866 -449 5888
rect -435 5894 -425 5903
rect -394 5896 -386 5903
rect -371 5895 -363 5929
rect -248 5903 -199 5911
rect -270 5866 -262 5888
rect -248 5894 -238 5903
rect -207 5896 -199 5903
rect -184 5895 -176 5929
rect -551 5853 -194 5854
rect -551 5845 -381 5853
rect -374 5846 -194 5853
rect -187 5846 -153 5854
rect -374 5845 -153 5846
rect -551 5843 -153 5845
rect -142 5835 -130 5929
rect -3 5929 125 5931
rect -67 5903 -18 5911
rect -89 5866 -81 5888
rect -67 5894 -57 5903
rect -26 5896 -18 5903
rect -3 5895 5 5929
rect 17 5928 125 5929
rect -142 5828 -13 5835
rect -6 5828 27 5835
rect -142 5825 27 5828
rect 103 5767 120 5928
rect 218 5789 237 6077
rect 1264 5818 1279 5819
rect 3207 5818 3215 5826
rect 1262 5809 3216 5818
rect 218 5788 343 5789
rect 1264 5788 1279 5809
rect 3207 5805 3215 5809
rect 218 5774 1280 5788
rect 103 5756 509 5767
rect 103 5754 518 5756
rect 1264 5763 1277 5774
rect 103 5753 338 5754
rect 1264 5753 1265 5763
rect 1276 5753 1277 5763
rect 766 5743 1025 5745
rect 489 5732 751 5742
rect 766 5736 1017 5743
rect 1024 5736 1025 5743
rect 1506 5737 1765 5739
rect 766 5735 1025 5736
rect -765 5701 -748 5710
rect 351 5709 398 5722
rect 501 5721 509 5732
rect 704 5721 712 5732
rect -765 5700 -709 5701
rect -765 5690 -702 5700
rect -1299 2459 -1297 2503
rect -1221 2500 -1216 2530
rect -1190 5679 -1172 5686
rect -899 5680 -857 5681
rect -944 5679 -827 5680
rect -1190 5671 -827 5679
rect -1190 5669 -925 5671
rect -899 5670 -857 5671
rect -1190 2495 -1172 5669
rect -765 5316 -749 5690
rect 386 5687 398 5709
rect 435 5715 509 5721
rect 435 5701 442 5715
rect 501 5699 509 5715
rect -710 5672 -703 5680
rect -300 5675 -41 5677
rect -656 5664 -315 5674
rect -300 5668 -49 5675
rect -42 5668 -41 5675
rect -300 5667 -41 5668
rect -565 5653 -557 5664
rect -362 5653 -354 5664
rect -631 5647 -557 5653
rect -631 5633 -624 5647
rect -565 5631 -557 5647
rect -428 5647 -354 5653
rect -428 5633 -421 5647
rect -609 5592 -600 5623
rect -362 5631 -354 5647
rect -546 5602 -538 5623
rect -547 5592 -538 5602
rect -609 5589 -538 5592
rect -406 5592 -397 5623
rect -343 5592 -335 5623
rect -406 5591 -335 5592
rect -299 5591 -290 5667
rect -175 5653 -167 5662
rect 6 5653 14 5662
rect -241 5647 -167 5653
rect -241 5633 -234 5647
rect -175 5631 -167 5647
rect -609 5584 -512 5589
rect -406 5584 -290 5591
rect -60 5647 14 5653
rect 389 5659 398 5687
rect 638 5715 712 5721
rect 638 5701 645 5715
rect 457 5660 466 5691
rect 704 5699 712 5715
rect 520 5670 528 5691
rect 519 5660 528 5670
rect 389 5656 453 5659
rect 389 5647 446 5656
rect -60 5633 -53 5647
rect -219 5592 -210 5623
rect 6 5631 14 5647
rect 457 5657 528 5660
rect 660 5660 669 5691
rect 723 5660 731 5691
rect 660 5659 731 5660
rect 767 5659 776 5735
rect 891 5721 899 5730
rect 1072 5721 1080 5730
rect 1150 5726 1491 5736
rect 1506 5730 1757 5737
rect 1764 5730 1765 5737
rect 1506 5729 1765 5730
rect 825 5715 899 5721
rect 825 5701 832 5715
rect 891 5699 899 5715
rect 457 5652 554 5657
rect 660 5652 776 5659
rect 1006 5715 1080 5721
rect 1241 5715 1249 5726
rect 1444 5715 1452 5726
rect 1006 5701 1013 5715
rect 847 5660 856 5691
rect 1072 5699 1080 5715
rect 910 5660 918 5691
rect 847 5659 918 5660
rect 1175 5709 1249 5715
rect 1028 5660 1037 5691
rect 1091 5660 1099 5691
rect 1175 5695 1182 5709
rect 1241 5693 1249 5709
rect 1028 5659 1099 5660
rect 1378 5709 1452 5715
rect 1378 5695 1385 5709
rect 847 5652 964 5659
rect 1028 5652 1122 5659
rect 520 5648 554 5652
rect -156 5592 -148 5623
rect -219 5591 -148 5592
rect -38 5592 -29 5623
rect 25 5592 33 5623
rect 456 5624 505 5632
rect -38 5591 33 5592
rect 41 5591 263 5594
rect -219 5584 -102 5591
rect -38 5584 263 5591
rect 434 5587 442 5609
rect 456 5615 466 5624
rect 497 5617 505 5624
rect 520 5616 528 5648
rect -546 5580 -512 5584
rect -610 5556 -561 5564
rect -632 5519 -624 5541
rect -610 5547 -600 5556
rect -569 5549 -561 5556
rect -546 5548 -538 5580
rect -523 5507 -512 5580
rect -343 5582 -290 5584
rect -156 5582 -102 5584
rect -407 5556 -358 5564
rect -429 5519 -421 5541
rect -407 5547 -397 5556
rect -366 5549 -358 5556
rect -343 5548 -335 5582
rect -220 5556 -171 5564
rect -242 5519 -234 5541
rect -220 5547 -210 5556
rect -179 5549 -171 5556
rect -156 5548 -148 5582
rect -523 5506 -166 5507
rect -523 5498 -353 5506
rect -346 5499 -166 5506
rect -159 5499 -125 5507
rect -346 5498 -125 5499
rect -523 5496 -125 5498
rect -114 5488 -102 5582
rect 25 5583 263 5584
rect 25 5582 53 5583
rect -39 5556 10 5564
rect -61 5519 -53 5541
rect -39 5547 -29 5556
rect 2 5549 10 5556
rect 25 5548 33 5582
rect -114 5481 15 5488
rect 22 5481 55 5488
rect -114 5478 55 5481
rect -768 5314 -715 5316
rect -768 5304 -702 5314
rect -768 5301 -715 5304
rect -1150 5284 -891 5295
rect -1150 2473 -1138 5284
rect -766 4891 -747 5301
rect -300 5289 -41 5291
rect -656 5278 -315 5288
rect -300 5282 -49 5289
rect -42 5282 -41 5289
rect -300 5281 -41 5282
rect -565 5267 -557 5278
rect -362 5267 -354 5278
rect -631 5261 -557 5267
rect -631 5247 -624 5261
rect -565 5245 -557 5261
rect -428 5261 -354 5267
rect -428 5247 -421 5261
rect -609 5206 -600 5237
rect -362 5245 -354 5261
rect -546 5216 -538 5237
rect -547 5206 -538 5216
rect -609 5203 -538 5206
rect -406 5206 -397 5237
rect -343 5206 -335 5237
rect -406 5205 -335 5206
rect -299 5205 -290 5281
rect -175 5267 -167 5276
rect 6 5267 14 5276
rect -241 5261 -167 5267
rect -241 5247 -234 5261
rect -175 5245 -167 5261
rect -609 5198 -512 5203
rect -406 5198 -290 5205
rect -60 5261 14 5267
rect -60 5247 -53 5261
rect -219 5206 -210 5237
rect 6 5245 14 5261
rect -156 5206 -148 5237
rect -219 5205 -148 5206
rect -38 5206 -29 5237
rect 25 5206 33 5237
rect -38 5205 33 5206
rect 92 5205 105 5206
rect -219 5198 -102 5205
rect -38 5198 109 5205
rect -546 5194 -512 5198
rect -610 5170 -561 5178
rect -632 5133 -624 5155
rect -610 5161 -600 5170
rect -569 5163 -561 5170
rect -546 5162 -538 5194
rect -523 5121 -512 5194
rect -343 5196 -290 5198
rect -156 5196 -102 5198
rect -407 5170 -358 5178
rect -429 5133 -421 5155
rect -407 5161 -397 5170
rect -366 5163 -358 5170
rect -343 5162 -335 5196
rect -220 5170 -171 5178
rect -242 5133 -234 5155
rect -220 5161 -210 5170
rect -179 5163 -171 5170
rect -156 5162 -148 5196
rect -523 5120 -166 5121
rect -523 5112 -353 5120
rect -346 5113 -166 5120
rect -159 5113 -125 5121
rect -346 5112 -125 5113
rect -523 5110 -125 5112
rect -114 5102 -102 5196
rect 25 5197 109 5198
rect 25 5196 53 5197
rect -39 5170 10 5178
rect -61 5133 -53 5155
rect -39 5161 -29 5170
rect 2 5163 10 5170
rect 25 5162 33 5196
rect -114 5095 15 5102
rect 22 5095 55 5102
rect -114 5092 55 5095
rect -766 4890 -713 4891
rect -766 4880 -702 4890
rect -766 4879 -713 4880
rect -735 4877 -713 4879
rect -1299 2458 -1274 2459
rect -1110 4870 -719 4871
rect -1110 4862 -703 4870
rect -300 4865 -41 4867
rect -1110 4861 -719 4862
rect -1110 2469 -1097 4861
rect -656 4854 -315 4864
rect -300 4858 -49 4865
rect -42 4858 -41 4865
rect -300 4857 -41 4858
rect -565 4843 -557 4854
rect -362 4843 -354 4854
rect -631 4837 -557 4843
rect -631 4823 -624 4837
rect -565 4821 -557 4837
rect -428 4837 -354 4843
rect -428 4823 -421 4837
rect -609 4782 -600 4813
rect -362 4821 -354 4837
rect -546 4792 -538 4813
rect -547 4782 -538 4792
rect -609 4779 -538 4782
rect -406 4782 -397 4813
rect -343 4782 -335 4813
rect -406 4781 -335 4782
rect -299 4781 -290 4857
rect -175 4843 -167 4852
rect 6 4843 14 4852
rect -241 4837 -167 4843
rect -241 4823 -234 4837
rect -175 4821 -167 4837
rect -609 4774 -512 4779
rect -406 4774 -290 4781
rect -60 4837 14 4843
rect -60 4823 -53 4837
rect -219 4782 -210 4813
rect 6 4821 14 4837
rect -156 4782 -148 4813
rect -219 4781 -148 4782
rect -38 4782 -29 4813
rect 25 4782 33 4813
rect -38 4781 33 4782
rect 44 4781 57 4783
rect -219 4774 -102 4781
rect -38 4774 57 4781
rect -546 4770 -512 4774
rect -610 4746 -561 4754
rect -632 4709 -624 4731
rect -610 4737 -600 4746
rect -569 4739 -561 4746
rect -546 4738 -538 4770
rect -523 4697 -512 4770
rect -343 4772 -290 4774
rect -156 4772 -102 4774
rect -407 4746 -358 4754
rect -429 4709 -421 4731
rect -407 4737 -397 4746
rect -366 4739 -358 4746
rect -343 4738 -335 4772
rect -220 4746 -171 4754
rect -242 4709 -234 4731
rect -220 4737 -210 4746
rect -179 4739 -171 4746
rect -156 4738 -148 4772
rect -523 4696 -166 4697
rect -523 4688 -353 4696
rect -346 4689 -166 4696
rect -159 4689 -125 4697
rect -346 4688 -125 4689
rect -523 4686 -125 4688
rect -114 4678 -102 4772
rect 25 4772 57 4774
rect -39 4746 10 4754
rect -61 4709 -53 4731
rect -39 4737 -29 4746
rect 2 4739 10 4746
rect 25 4738 33 4772
rect -114 4671 15 4678
rect 22 4671 30 4678
rect -114 4668 30 4671
rect 44 3831 57 4772
rect 92 4405 105 5197
rect 245 5044 262 5583
rect 543 5575 554 5648
rect 723 5650 776 5652
rect 910 5650 964 5652
rect 659 5624 708 5632
rect 637 5587 645 5609
rect 659 5615 669 5624
rect 700 5617 708 5624
rect 723 5616 731 5650
rect 846 5624 895 5632
rect 824 5587 832 5609
rect 846 5615 856 5624
rect 887 5617 895 5624
rect 910 5616 918 5650
rect 543 5574 900 5575
rect 543 5566 713 5574
rect 720 5567 900 5574
rect 907 5567 941 5575
rect 720 5566 941 5567
rect 543 5564 941 5566
rect 952 5556 964 5650
rect 1091 5650 1122 5652
rect 1027 5624 1076 5632
rect 1005 5587 1013 5609
rect 1027 5615 1037 5624
rect 1068 5617 1076 5624
rect 1091 5616 1099 5650
rect 1114 5644 1122 5650
rect 1197 5654 1206 5685
rect 1444 5693 1452 5709
rect 1260 5664 1268 5685
rect 1259 5654 1268 5664
rect 1197 5651 1268 5654
rect 1400 5654 1409 5685
rect 1463 5654 1471 5685
rect 1400 5653 1471 5654
rect 1507 5653 1516 5729
rect 1631 5715 1639 5724
rect 1812 5715 1820 5724
rect 1565 5709 1639 5715
rect 1565 5695 1572 5709
rect 1631 5693 1639 5709
rect 1197 5646 1294 5651
rect 1400 5646 1516 5653
rect 1746 5709 1820 5715
rect 2257 5713 2265 5718
rect 1746 5695 1753 5709
rect 1587 5654 1596 5685
rect 1812 5693 1820 5709
rect 1650 5654 1658 5685
rect 1587 5653 1658 5654
rect 2191 5707 2265 5713
rect 2191 5693 2198 5707
rect 1768 5654 1777 5685
rect 2257 5691 2265 5707
rect 2397 5703 2405 5711
rect 3033 5704 3040 5720
rect 1831 5654 1839 5685
rect 1768 5653 1839 5654
rect 2362 5697 2405 5703
rect 1587 5646 1704 5653
rect 1768 5646 2202 5653
rect 1114 5636 1185 5644
rect 1114 5635 1194 5636
rect 1260 5642 1294 5646
rect 952 5549 1081 5556
rect 1088 5549 1121 5556
rect 952 5546 1121 5549
rect 1136 5528 1149 5635
rect 1196 5618 1245 5626
rect 1174 5581 1182 5603
rect 1196 5609 1206 5618
rect 1237 5611 1245 5618
rect 1260 5610 1268 5642
rect 1283 5569 1294 5642
rect 1463 5644 1516 5646
rect 1650 5644 1704 5646
rect 1399 5618 1448 5626
rect 1377 5581 1385 5603
rect 1399 5609 1409 5618
rect 1440 5611 1448 5618
rect 1463 5610 1471 5644
rect 1586 5618 1635 5626
rect 1564 5581 1572 5603
rect 1586 5609 1596 5618
rect 1627 5611 1635 5618
rect 1650 5610 1658 5644
rect 1283 5568 1640 5569
rect 1283 5560 1453 5568
rect 1460 5561 1640 5568
rect 1647 5561 1681 5569
rect 1460 5560 1681 5561
rect 1283 5558 1681 5560
rect 1692 5550 1704 5644
rect 1831 5645 2202 5646
rect 2209 5645 2210 5653
rect 2213 5652 2222 5683
rect 2362 5683 2370 5697
rect 2276 5652 2284 5683
rect 2213 5650 2284 5652
rect 3050 5674 3058 5695
rect 3158 5674 3165 5752
rect 3204 5691 3218 5805
rect 3277 5691 3288 5693
rect 3204 5677 3288 5691
rect 2213 5649 2285 5650
rect 1831 5644 1850 5645
rect 2017 5644 2036 5645
rect 2213 5644 2310 5649
rect 1767 5618 1816 5626
rect 1745 5581 1753 5603
rect 1767 5609 1777 5618
rect 1808 5611 1816 5618
rect 1831 5610 1839 5644
rect 2276 5640 2310 5644
rect 2212 5616 2261 5624
rect 1879 5610 2037 5613
rect 1878 5599 2037 5610
rect 1878 5597 1901 5599
rect 1957 5597 2037 5599
rect 1692 5543 1821 5550
rect 1828 5543 1861 5550
rect 1692 5540 1861 5543
rect 455 5516 1152 5528
rect 458 5503 468 5516
rect 1878 5511 1894 5597
rect 2190 5579 2198 5601
rect 2212 5607 2222 5616
rect 2253 5609 2261 5616
rect 2276 5608 2284 5640
rect 2299 5635 2310 5640
rect 2385 5637 2395 5670
rect 2299 5625 2340 5635
rect 2385 5628 2990 5637
rect 2385 5602 2395 5628
rect 2361 5575 2370 5591
rect 2361 5569 2396 5575
rect 456 5487 468 5503
rect 1793 5498 1934 5511
rect 456 5473 457 5487
rect 467 5473 468 5487
rect 401 5429 409 5434
rect 335 5423 409 5429
rect 335 5409 342 5423
rect 401 5407 409 5423
rect 541 5419 549 5427
rect 506 5413 549 5419
rect 584 5415 593 5478
rect 749 5439 756 5473
rect 700 5433 756 5439
rect 684 5425 692 5430
rect 357 5368 366 5399
rect 506 5399 514 5413
rect 618 5419 692 5425
rect 618 5405 625 5419
rect 684 5403 692 5419
rect 824 5415 832 5423
rect 420 5368 428 5399
rect 357 5366 428 5368
rect 357 5365 429 5366
rect 357 5360 454 5365
rect 420 5356 454 5360
rect 356 5332 405 5340
rect 334 5295 342 5317
rect 356 5323 366 5332
rect 397 5325 405 5332
rect 420 5324 428 5356
rect 443 5351 454 5356
rect 529 5353 539 5386
rect 789 5409 832 5415
rect 640 5364 649 5395
rect 789 5395 797 5409
rect 880 5407 903 5413
rect 880 5397 886 5407
rect 703 5364 711 5395
rect 640 5362 711 5364
rect 971 5397 977 5413
rect 640 5361 712 5362
rect 640 5356 737 5361
rect 443 5341 484 5351
rect 529 5344 546 5353
rect 529 5318 539 5344
rect 554 5344 556 5353
rect 703 5352 737 5356
rect 639 5328 688 5336
rect 505 5291 514 5307
rect 617 5291 625 5313
rect 639 5319 649 5328
rect 680 5321 688 5328
rect 703 5320 711 5352
rect 726 5347 737 5352
rect 812 5349 822 5382
rect 899 5375 905 5388
rect 920 5375 926 5388
rect 899 5369 926 5375
rect 940 5366 946 5388
rect 989 5368 996 5389
rect 1793 5368 1802 5498
rect 940 5360 962 5366
rect 989 5360 1802 5368
rect 940 5354 946 5360
rect 726 5337 767 5347
rect 812 5341 850 5349
rect 899 5348 946 5354
rect 812 5340 849 5341
rect 812 5314 822 5340
rect 505 5285 540 5291
rect 788 5287 797 5303
rect 788 5281 823 5287
rect 838 5251 849 5340
rect 899 5336 906 5348
rect 939 5336 946 5348
rect 989 5359 1793 5360
rect 989 5336 996 5359
rect 880 5316 886 5330
rect 920 5316 926 5330
rect 880 5311 949 5316
rect 971 5313 977 5330
rect 1066 5064 1089 5359
rect 391 5050 1337 5064
rect 243 5043 404 5044
rect 243 5032 566 5043
rect 243 5030 575 5032
rect 1321 5039 1334 5050
rect 327 5029 404 5030
rect 1321 5029 1322 5039
rect 1333 5029 1334 5039
rect 823 5019 1082 5021
rect 546 5008 808 5018
rect 823 5012 1074 5019
rect 1081 5012 1082 5019
rect 1563 5013 1822 5015
rect 823 5011 1082 5012
rect 409 4985 455 4998
rect 558 4997 566 5008
rect 761 4997 769 5008
rect 443 4963 455 4985
rect 492 4991 566 4997
rect 492 4977 499 4991
rect 558 4975 566 4991
rect 446 4935 455 4963
rect 695 4991 769 4997
rect 695 4977 702 4991
rect 514 4936 523 4967
rect 761 4975 769 4991
rect 577 4946 585 4967
rect 576 4936 585 4946
rect 446 4932 510 4935
rect 446 4923 503 4932
rect 514 4933 585 4936
rect 717 4936 726 4967
rect 780 4936 788 4967
rect 717 4935 788 4936
rect 824 4935 833 5011
rect 948 4997 956 5006
rect 1129 4997 1137 5006
rect 1207 5002 1548 5012
rect 1563 5006 1814 5013
rect 1821 5006 1822 5013
rect 1563 5005 1822 5006
rect 882 4991 956 4997
rect 882 4977 889 4991
rect 948 4975 956 4991
rect 514 4928 611 4933
rect 717 4928 833 4935
rect 1063 4991 1137 4997
rect 1298 4991 1306 5002
rect 1501 4991 1509 5002
rect 1063 4977 1070 4991
rect 904 4936 913 4967
rect 1129 4975 1137 4991
rect 967 4936 975 4967
rect 904 4935 975 4936
rect 1232 4985 1306 4991
rect 1085 4936 1094 4967
rect 1148 4936 1156 4967
rect 1232 4971 1239 4985
rect 1298 4969 1306 4985
rect 1085 4935 1156 4936
rect 1435 4985 1509 4991
rect 1435 4971 1442 4985
rect 904 4928 1021 4935
rect 1085 4928 1179 4935
rect 577 4924 611 4928
rect 513 4900 562 4908
rect 491 4863 499 4885
rect 513 4891 523 4900
rect 554 4893 562 4900
rect 577 4892 585 4924
rect 600 4851 611 4924
rect 780 4926 833 4928
rect 967 4926 1021 4928
rect 716 4900 765 4908
rect 694 4863 702 4885
rect 716 4891 726 4900
rect 757 4893 765 4900
rect 780 4892 788 4926
rect 903 4900 952 4908
rect 881 4863 889 4885
rect 903 4891 913 4900
rect 944 4893 952 4900
rect 967 4892 975 4926
rect 600 4850 957 4851
rect 600 4842 770 4850
rect 777 4843 957 4850
rect 964 4843 998 4851
rect 777 4842 998 4843
rect 600 4840 998 4842
rect 1009 4832 1021 4926
rect 1148 4926 1179 4928
rect 1084 4900 1133 4908
rect 1062 4863 1070 4885
rect 1084 4891 1094 4900
rect 1125 4893 1133 4900
rect 1148 4892 1156 4926
rect 1171 4920 1179 4926
rect 1254 4930 1263 4961
rect 1501 4969 1509 4985
rect 1317 4940 1325 4961
rect 1316 4930 1325 4940
rect 1254 4927 1325 4930
rect 1457 4930 1466 4961
rect 1520 4930 1528 4961
rect 1457 4929 1528 4930
rect 1564 4929 1573 5005
rect 1688 4991 1696 5000
rect 1869 4991 1877 5000
rect 1622 4985 1696 4991
rect 1622 4971 1629 4985
rect 1688 4969 1696 4985
rect 1254 4922 1351 4927
rect 1457 4922 1573 4929
rect 1803 4985 1877 4991
rect 2255 4989 2263 4994
rect 1803 4971 1810 4985
rect 1644 4930 1653 4961
rect 1869 4969 1877 4985
rect 1707 4930 1715 4961
rect 1644 4929 1715 4930
rect 2189 4983 2263 4989
rect 2189 4969 2196 4983
rect 1825 4930 1834 4961
rect 2255 4967 2263 4983
rect 2395 4979 2403 4987
rect 1888 4930 1896 4961
rect 2360 4973 2403 4979
rect 1825 4929 1896 4930
rect 1994 4929 2145 4930
rect 1644 4922 1761 4929
rect 1825 4922 2200 4929
rect 1171 4912 1242 4920
rect 1171 4911 1251 4912
rect 1317 4918 1351 4922
rect 1009 4825 1138 4832
rect 1145 4825 1178 4832
rect 1009 4822 1178 4825
rect 1193 4804 1206 4911
rect 1253 4894 1302 4902
rect 1231 4857 1239 4879
rect 1253 4885 1263 4894
rect 1294 4887 1302 4894
rect 1317 4886 1325 4918
rect 1340 4845 1351 4918
rect 1520 4920 1573 4922
rect 1707 4920 1761 4922
rect 1456 4894 1505 4902
rect 1434 4857 1442 4879
rect 1456 4885 1466 4894
rect 1497 4887 1505 4894
rect 1520 4886 1528 4920
rect 1643 4894 1692 4902
rect 1621 4857 1629 4879
rect 1643 4885 1653 4894
rect 1684 4887 1692 4894
rect 1707 4886 1715 4920
rect 1340 4844 1697 4845
rect 1340 4836 1510 4844
rect 1517 4837 1697 4844
rect 1704 4837 1738 4845
rect 1517 4836 1738 4837
rect 1340 4834 1738 4836
rect 1749 4826 1761 4920
rect 1888 4921 2200 4922
rect 2207 4921 2208 4929
rect 2211 4928 2220 4959
rect 2360 4959 2368 4973
rect 2274 4928 2282 4959
rect 2211 4926 2282 4928
rect 2211 4925 2283 4926
rect 1888 4920 1907 4921
rect 2211 4920 2308 4925
rect 1824 4894 1873 4902
rect 1802 4857 1810 4879
rect 1824 4885 1834 4894
rect 1865 4887 1873 4894
rect 1888 4886 1896 4920
rect 2274 4916 2308 4920
rect 2210 4892 2259 4900
rect 1936 4886 2094 4889
rect 1935 4875 2094 4886
rect 1935 4873 1958 4875
rect 2014 4873 2094 4875
rect 1749 4819 1878 4826
rect 1885 4819 1918 4826
rect 1749 4816 1918 4819
rect 512 4792 1209 4804
rect 515 4779 525 4792
rect 1935 4787 1951 4873
rect 2188 4855 2196 4877
rect 2210 4883 2220 4892
rect 2251 4885 2259 4892
rect 2274 4884 2282 4916
rect 2297 4911 2308 4916
rect 2383 4913 2393 4946
rect 2383 4912 2786 4913
rect 2297 4901 2338 4911
rect 2383 4904 2946 4912
rect 2383 4878 2393 4904
rect 2403 4903 2946 4904
rect 2403 4902 2786 4903
rect 2359 4851 2368 4867
rect 2359 4845 2394 4851
rect 513 4763 525 4779
rect 1850 4774 1991 4787
rect 513 4749 514 4763
rect 524 4749 525 4763
rect 458 4705 466 4710
rect 392 4699 466 4705
rect 392 4685 399 4699
rect 458 4683 466 4699
rect 598 4695 606 4703
rect 563 4689 606 4695
rect 641 4691 650 4754
rect 806 4715 813 4749
rect 757 4709 813 4715
rect 741 4701 749 4706
rect 414 4644 423 4675
rect 563 4675 571 4689
rect 675 4695 749 4701
rect 675 4681 682 4695
rect 741 4679 749 4695
rect 881 4691 889 4699
rect 477 4644 485 4675
rect 414 4642 485 4644
rect 414 4641 486 4642
rect 414 4636 511 4641
rect 477 4632 511 4636
rect 413 4608 462 4616
rect 391 4571 399 4593
rect 413 4599 423 4608
rect 454 4601 462 4608
rect 477 4600 485 4632
rect 500 4627 511 4632
rect 586 4629 596 4662
rect 846 4685 889 4691
rect 697 4640 706 4671
rect 846 4671 854 4685
rect 937 4683 960 4689
rect 937 4673 943 4683
rect 760 4640 768 4671
rect 697 4638 768 4640
rect 1028 4673 1034 4689
rect 697 4637 769 4638
rect 697 4632 794 4637
rect 500 4617 541 4627
rect 586 4620 603 4629
rect 586 4594 596 4620
rect 611 4620 613 4629
rect 760 4628 794 4632
rect 696 4604 745 4612
rect 562 4567 571 4583
rect 674 4567 682 4589
rect 696 4595 706 4604
rect 737 4597 745 4604
rect 760 4596 768 4628
rect 783 4623 794 4628
rect 869 4625 879 4658
rect 956 4651 962 4664
rect 977 4651 983 4664
rect 956 4645 983 4651
rect 997 4642 1003 4664
rect 1046 4644 1053 4665
rect 1850 4644 1859 4774
rect 997 4636 1019 4642
rect 1046 4636 1859 4644
rect 997 4630 1003 4636
rect 783 4613 824 4623
rect 869 4617 907 4625
rect 956 4624 1003 4630
rect 869 4616 906 4617
rect 869 4590 879 4616
rect 562 4561 597 4567
rect 845 4563 854 4579
rect 845 4557 880 4563
rect 895 4527 906 4616
rect 956 4612 963 4624
rect 996 4612 1003 4624
rect 1046 4635 1850 4636
rect 1046 4612 1053 4635
rect 937 4592 943 4606
rect 977 4592 983 4606
rect 937 4587 1006 4592
rect 1028 4589 1034 4606
rect 1154 4474 1167 4635
rect 371 4460 1317 4474
rect 134 4453 387 4454
rect 134 4442 546 4453
rect 134 4440 555 4442
rect 1301 4449 1314 4460
rect 134 4437 387 4440
rect 1301 4439 1302 4449
rect 1313 4439 1314 4449
rect 803 4429 1062 4431
rect 526 4418 788 4428
rect 803 4422 1054 4429
rect 1061 4422 1062 4429
rect 1543 4423 1802 4425
rect 803 4421 1062 4422
rect 371 4405 435 4408
rect 538 4407 546 4418
rect 741 4407 749 4418
rect 92 4396 435 4405
rect 92 4395 381 4396
rect 388 4395 435 4396
rect 92 4386 105 4395
rect 423 4373 435 4395
rect 472 4401 546 4407
rect 472 4387 479 4401
rect 538 4385 546 4401
rect 426 4345 435 4373
rect 675 4401 749 4407
rect 675 4387 682 4401
rect 494 4346 503 4377
rect 741 4385 749 4401
rect 557 4356 565 4377
rect 556 4346 565 4356
rect 426 4342 490 4345
rect 426 4333 483 4342
rect 494 4343 565 4346
rect 697 4346 706 4377
rect 760 4346 768 4377
rect 697 4345 768 4346
rect 804 4345 813 4421
rect 928 4407 936 4416
rect 1109 4407 1117 4416
rect 1187 4412 1528 4422
rect 1543 4416 1794 4423
rect 1801 4416 1802 4423
rect 1543 4415 1802 4416
rect 862 4401 936 4407
rect 862 4387 869 4401
rect 928 4385 936 4401
rect 494 4338 591 4343
rect 697 4338 813 4345
rect 1043 4401 1117 4407
rect 1278 4401 1286 4412
rect 1481 4401 1489 4412
rect 1043 4387 1050 4401
rect 884 4346 893 4377
rect 1109 4385 1117 4401
rect 947 4346 955 4377
rect 884 4345 955 4346
rect 1212 4395 1286 4401
rect 1065 4346 1074 4377
rect 1128 4346 1136 4377
rect 1212 4381 1219 4395
rect 1278 4379 1286 4395
rect 1065 4345 1136 4346
rect 1415 4395 1489 4401
rect 1415 4381 1422 4395
rect 884 4338 1001 4345
rect 1065 4338 1159 4345
rect 557 4334 591 4338
rect 493 4310 542 4318
rect 471 4273 479 4295
rect 493 4301 503 4310
rect 534 4303 542 4310
rect 557 4302 565 4334
rect 580 4261 591 4334
rect 760 4336 813 4338
rect 947 4336 1001 4338
rect 696 4310 745 4318
rect 674 4273 682 4295
rect 696 4301 706 4310
rect 737 4303 745 4310
rect 760 4302 768 4336
rect 883 4310 932 4318
rect 861 4273 869 4295
rect 883 4301 893 4310
rect 924 4303 932 4310
rect 947 4302 955 4336
rect 580 4260 937 4261
rect 580 4252 750 4260
rect 757 4253 937 4260
rect 944 4253 978 4261
rect 757 4252 978 4253
rect 580 4250 978 4252
rect 989 4242 1001 4336
rect 1128 4336 1159 4338
rect 1064 4310 1113 4318
rect 1042 4273 1050 4295
rect 1064 4301 1074 4310
rect 1105 4303 1113 4310
rect 1128 4302 1136 4336
rect 1151 4330 1159 4336
rect 1234 4340 1243 4371
rect 1481 4379 1489 4395
rect 1297 4350 1305 4371
rect 1296 4340 1305 4350
rect 1234 4337 1305 4340
rect 1437 4340 1446 4371
rect 1500 4340 1508 4371
rect 1437 4339 1508 4340
rect 1544 4339 1553 4415
rect 1668 4401 1676 4410
rect 1849 4401 1857 4410
rect 1602 4395 1676 4401
rect 1602 4381 1609 4395
rect 1668 4379 1676 4395
rect 1234 4332 1331 4337
rect 1437 4332 1553 4339
rect 1783 4395 1857 4401
rect 2256 4399 2264 4404
rect 1783 4381 1790 4395
rect 1624 4340 1633 4371
rect 1849 4379 1857 4395
rect 1687 4340 1695 4371
rect 1624 4339 1695 4340
rect 2190 4393 2264 4399
rect 2190 4379 2197 4393
rect 1805 4340 1814 4371
rect 2256 4377 2264 4393
rect 2396 4389 2404 4397
rect 1868 4340 1876 4371
rect 2361 4383 2404 4389
rect 1805 4339 1876 4340
rect 2055 4339 2146 4340
rect 1624 4332 1741 4339
rect 1805 4332 2201 4339
rect 1151 4322 1222 4330
rect 1151 4321 1231 4322
rect 1297 4328 1331 4332
rect 989 4235 1118 4242
rect 1125 4235 1158 4242
rect 989 4232 1158 4235
rect 1173 4214 1186 4321
rect 1233 4304 1282 4312
rect 1211 4267 1219 4289
rect 1233 4295 1243 4304
rect 1274 4297 1282 4304
rect 1297 4296 1305 4328
rect 1320 4255 1331 4328
rect 1500 4330 1553 4332
rect 1687 4330 1741 4332
rect 1436 4304 1485 4312
rect 1414 4267 1422 4289
rect 1436 4295 1446 4304
rect 1477 4297 1485 4304
rect 1500 4296 1508 4330
rect 1623 4304 1672 4312
rect 1601 4267 1609 4289
rect 1623 4295 1633 4304
rect 1664 4297 1672 4304
rect 1687 4296 1695 4330
rect 1320 4254 1677 4255
rect 1320 4246 1490 4254
rect 1497 4247 1677 4254
rect 1684 4247 1718 4255
rect 1497 4246 1718 4247
rect 1320 4244 1718 4246
rect 1729 4236 1741 4330
rect 1868 4331 2201 4332
rect 2208 4331 2209 4339
rect 2212 4338 2221 4369
rect 2361 4369 2369 4383
rect 2275 4338 2283 4369
rect 2212 4336 2283 4338
rect 2212 4335 2284 4336
rect 1868 4330 1887 4331
rect 2212 4330 2309 4335
rect 1804 4304 1853 4312
rect 1782 4267 1790 4289
rect 1804 4295 1814 4304
rect 1845 4297 1853 4304
rect 1868 4296 1876 4330
rect 2275 4326 2309 4330
rect 2211 4302 2260 4310
rect 2046 4299 2074 4300
rect 1916 4296 2074 4299
rect 1915 4285 2074 4296
rect 1915 4283 1938 4285
rect 1994 4283 2074 4285
rect 1729 4229 1858 4236
rect 1865 4229 1898 4236
rect 1729 4226 1898 4229
rect 492 4202 1189 4214
rect 495 4189 505 4202
rect 1915 4197 1931 4283
rect 2189 4265 2197 4287
rect 2211 4293 2221 4302
rect 2252 4295 2260 4302
rect 2275 4294 2283 4326
rect 2298 4321 2309 4326
rect 2384 4323 2394 4356
rect 2444 4324 2727 4325
rect 2409 4323 2887 4324
rect 2298 4311 2339 4321
rect 2384 4315 2887 4323
rect 2384 4314 2727 4315
rect 2384 4288 2394 4314
rect 2409 4313 2481 4314
rect 2360 4261 2369 4277
rect 2360 4255 2395 4261
rect 493 4173 505 4189
rect 1830 4184 1971 4197
rect 493 4159 494 4173
rect 504 4159 505 4173
rect 438 4115 446 4120
rect 372 4109 446 4115
rect 372 4095 379 4109
rect 438 4093 446 4109
rect 578 4105 586 4113
rect 543 4099 586 4105
rect 621 4101 630 4164
rect 786 4125 793 4159
rect 737 4119 793 4125
rect 721 4111 729 4116
rect 394 4054 403 4085
rect 543 4085 551 4099
rect 655 4105 729 4111
rect 655 4091 662 4105
rect 721 4089 729 4105
rect 861 4101 869 4109
rect 457 4054 465 4085
rect 394 4052 465 4054
rect 394 4051 466 4052
rect 394 4046 491 4051
rect 457 4042 491 4046
rect 393 4018 442 4026
rect 371 3981 379 4003
rect 393 4009 403 4018
rect 434 4011 442 4018
rect 457 4010 465 4042
rect 480 4037 491 4042
rect 566 4039 576 4072
rect 826 4095 869 4101
rect 677 4050 686 4081
rect 826 4081 834 4095
rect 917 4093 940 4099
rect 917 4083 923 4093
rect 740 4050 748 4081
rect 677 4048 748 4050
rect 1008 4083 1014 4099
rect 677 4047 749 4048
rect 677 4042 774 4047
rect 480 4027 521 4037
rect 566 4030 583 4039
rect 566 4004 576 4030
rect 591 4030 593 4039
rect 740 4038 774 4042
rect 676 4014 725 4022
rect 542 3977 551 3993
rect 654 3977 662 3999
rect 676 4005 686 4014
rect 717 4007 725 4014
rect 740 4006 748 4038
rect 763 4033 774 4038
rect 849 4035 859 4068
rect 936 4061 942 4074
rect 957 4061 963 4074
rect 936 4055 963 4061
rect 977 4052 983 4074
rect 1026 4054 1033 4075
rect 1830 4054 1839 4184
rect 977 4046 999 4052
rect 1026 4046 1839 4054
rect 977 4040 983 4046
rect 763 4023 804 4033
rect 849 4027 887 4035
rect 936 4034 983 4040
rect 849 4026 886 4027
rect 849 4000 859 4026
rect 542 3971 577 3977
rect 825 3973 834 3989
rect 825 3967 860 3973
rect 875 3937 886 4026
rect 936 4022 943 4034
rect 976 4022 983 4034
rect 1026 4045 1830 4046
rect 1026 4022 1033 4045
rect 917 4002 923 4016
rect 957 4002 963 4016
rect 917 3997 986 4002
rect 1008 3999 1014 4016
rect 1194 3850 1208 4045
rect 399 3836 1345 3850
rect 41 3829 411 3831
rect 41 3818 574 3829
rect 41 3816 583 3818
rect 1329 3825 1342 3836
rect 41 3815 411 3816
rect 1329 3815 1330 3825
rect 1341 3815 1342 3825
rect 831 3805 1090 3807
rect 554 3794 816 3804
rect 831 3798 1082 3805
rect 1089 3798 1090 3805
rect 1571 3799 1830 3801
rect 831 3797 1090 3798
rect 61 3784 402 3785
rect 61 3771 74 3784
rect 85 3772 463 3784
rect 566 3783 574 3794
rect 769 3783 777 3794
rect 85 3771 402 3772
rect 416 3771 463 3772
rect 451 3749 463 3771
rect 500 3777 574 3783
rect 500 3763 507 3777
rect 566 3761 574 3777
rect 454 3721 463 3749
rect 703 3777 777 3783
rect 703 3763 710 3777
rect 522 3722 531 3753
rect 769 3761 777 3777
rect 585 3732 593 3753
rect 584 3722 593 3732
rect 454 3718 518 3721
rect 454 3709 511 3718
rect 522 3719 593 3722
rect 725 3722 734 3753
rect 788 3722 796 3753
rect 725 3721 796 3722
rect 832 3721 841 3797
rect 956 3783 964 3792
rect 1137 3783 1145 3792
rect 1215 3788 1556 3798
rect 1571 3792 1822 3799
rect 1829 3792 1830 3799
rect 1571 3791 1830 3792
rect 890 3777 964 3783
rect 890 3763 897 3777
rect 956 3761 964 3777
rect 522 3714 619 3719
rect 725 3714 841 3721
rect 1071 3777 1145 3783
rect 1306 3777 1314 3788
rect 1509 3777 1517 3788
rect 1071 3763 1078 3777
rect 912 3722 921 3753
rect 1137 3761 1145 3777
rect 975 3722 983 3753
rect 912 3721 983 3722
rect 1240 3771 1314 3777
rect 1093 3722 1102 3753
rect 1156 3722 1164 3753
rect 1240 3757 1247 3771
rect 1306 3755 1314 3771
rect 1093 3721 1164 3722
rect 1443 3771 1517 3777
rect 1443 3757 1450 3771
rect 912 3714 1029 3721
rect 1093 3714 1187 3721
rect 585 3710 619 3714
rect 521 3686 570 3694
rect 499 3649 507 3671
rect 521 3677 531 3686
rect 562 3679 570 3686
rect 585 3678 593 3710
rect 608 3637 619 3710
rect 788 3712 841 3714
rect 975 3712 1029 3714
rect 724 3686 773 3694
rect 702 3649 710 3671
rect 724 3677 734 3686
rect 765 3679 773 3686
rect 788 3678 796 3712
rect 911 3686 960 3694
rect 889 3649 897 3671
rect 911 3677 921 3686
rect 952 3679 960 3686
rect 975 3678 983 3712
rect 608 3636 965 3637
rect 608 3628 778 3636
rect 785 3629 965 3636
rect 972 3629 1006 3637
rect 785 3628 1006 3629
rect 608 3626 1006 3628
rect 1017 3618 1029 3712
rect 1156 3712 1187 3714
rect 1092 3686 1141 3694
rect 1070 3649 1078 3671
rect 1092 3677 1102 3686
rect 1133 3679 1141 3686
rect 1156 3678 1164 3712
rect 1179 3706 1187 3712
rect 1262 3716 1271 3747
rect 1509 3755 1517 3771
rect 1325 3726 1333 3747
rect 1324 3716 1333 3726
rect 1262 3713 1333 3716
rect 1465 3716 1474 3747
rect 1528 3716 1536 3747
rect 1465 3715 1536 3716
rect 1572 3715 1581 3791
rect 1696 3777 1704 3786
rect 1877 3777 1885 3786
rect 1630 3771 1704 3777
rect 1630 3757 1637 3771
rect 1696 3755 1704 3771
rect 1262 3708 1359 3713
rect 1465 3708 1581 3715
rect 1811 3771 1885 3777
rect 2257 3775 2265 3780
rect 1811 3757 1818 3771
rect 1652 3716 1661 3747
rect 1877 3755 1885 3771
rect 1715 3716 1723 3747
rect 1652 3715 1723 3716
rect 2191 3769 2265 3775
rect 2191 3755 2198 3769
rect 1833 3716 1842 3747
rect 2257 3753 2265 3769
rect 2397 3765 2405 3773
rect 1896 3716 1904 3747
rect 1833 3715 1904 3716
rect 2362 3759 2405 3765
rect 1652 3708 1769 3715
rect 1833 3708 2202 3715
rect 1179 3698 1250 3706
rect 1179 3697 1259 3698
rect 1325 3704 1359 3708
rect 1017 3611 1146 3618
rect 1153 3611 1186 3618
rect 1017 3608 1186 3611
rect 1201 3590 1214 3697
rect 1261 3680 1310 3688
rect 1239 3643 1247 3665
rect 1261 3671 1271 3680
rect 1302 3673 1310 3680
rect 1325 3672 1333 3704
rect 1348 3631 1359 3704
rect 1528 3706 1581 3708
rect 1715 3706 1769 3708
rect 1464 3680 1513 3688
rect 1442 3643 1450 3665
rect 1464 3671 1474 3680
rect 1505 3673 1513 3680
rect 1528 3672 1536 3706
rect 1651 3680 1700 3688
rect 1629 3643 1637 3665
rect 1651 3671 1661 3680
rect 1692 3673 1700 3680
rect 1715 3672 1723 3706
rect 1348 3630 1705 3631
rect 1348 3622 1518 3630
rect 1525 3623 1705 3630
rect 1712 3623 1746 3631
rect 1525 3622 1746 3623
rect 1348 3620 1746 3622
rect 1757 3612 1769 3706
rect 1896 3707 2202 3708
rect 2209 3707 2210 3715
rect 2213 3714 2222 3745
rect 2362 3745 2370 3759
rect 2276 3714 2284 3745
rect 2213 3712 2284 3714
rect 2213 3711 2285 3712
rect 1896 3706 1915 3707
rect 2213 3706 2310 3711
rect 1832 3680 1881 3688
rect 1810 3643 1818 3665
rect 1832 3671 1842 3680
rect 1873 3673 1881 3680
rect 1896 3672 1904 3706
rect 2276 3702 2310 3706
rect 2212 3678 2261 3686
rect 1944 3672 2109 3675
rect 1943 3661 2109 3672
rect 1943 3659 1966 3661
rect 2022 3659 2109 3661
rect 1757 3605 1886 3612
rect 1893 3605 1926 3612
rect 1757 3602 1926 3605
rect 520 3578 1217 3590
rect 523 3565 533 3578
rect 1943 3573 1959 3659
rect 521 3549 533 3565
rect 1858 3560 1999 3573
rect 521 3535 522 3549
rect 532 3535 533 3549
rect 466 3491 474 3496
rect 400 3485 474 3491
rect 400 3471 407 3485
rect 466 3469 474 3485
rect 606 3481 614 3489
rect 571 3475 614 3481
rect 649 3477 658 3540
rect 814 3501 821 3535
rect 765 3495 821 3501
rect 749 3487 757 3492
rect 422 3430 431 3461
rect 571 3461 579 3475
rect 683 3481 757 3487
rect 683 3467 690 3481
rect 749 3465 757 3481
rect 889 3477 897 3485
rect 485 3430 493 3461
rect 422 3428 493 3430
rect 422 3427 494 3428
rect 422 3422 519 3427
rect 485 3418 519 3422
rect 421 3394 470 3402
rect 399 3357 407 3379
rect 421 3385 431 3394
rect 462 3387 470 3394
rect 485 3386 493 3418
rect 508 3413 519 3418
rect 594 3415 604 3448
rect 854 3471 897 3477
rect 705 3426 714 3457
rect 854 3457 862 3471
rect 945 3469 968 3475
rect 945 3459 951 3469
rect 768 3426 776 3457
rect 705 3424 776 3426
rect 1036 3459 1042 3475
rect 705 3423 777 3424
rect 705 3418 802 3423
rect 508 3403 549 3413
rect 594 3406 611 3415
rect 594 3380 604 3406
rect 619 3406 621 3415
rect 768 3414 802 3418
rect 704 3390 753 3398
rect 570 3353 579 3369
rect 682 3353 690 3375
rect 704 3381 714 3390
rect 745 3383 753 3390
rect 768 3382 776 3414
rect 791 3409 802 3414
rect 877 3411 887 3444
rect 964 3437 970 3450
rect 985 3437 991 3450
rect 964 3431 991 3437
rect 1005 3428 1011 3450
rect 1054 3430 1061 3451
rect 1858 3430 1867 3560
rect 2098 3539 2109 3659
rect 2190 3641 2198 3663
rect 2212 3669 2222 3678
rect 2253 3671 2261 3678
rect 2276 3670 2284 3702
rect 2299 3697 2310 3702
rect 2385 3699 2395 3732
rect 2299 3687 2340 3697
rect 2385 3690 2405 3699
rect 2385 3664 2395 3690
rect 2361 3637 2370 3653
rect 2361 3631 2396 3637
rect 2259 3599 2267 3604
rect 2193 3593 2267 3599
rect 2869 3601 2879 4315
rect 2928 4189 2938 4903
rect 2193 3579 2200 3593
rect 2259 3577 2267 3593
rect 2399 3589 2407 3597
rect 2364 3583 2407 3589
rect 2098 3531 2204 3539
rect 2211 3531 2212 3539
rect 2215 3538 2224 3569
rect 2364 3569 2372 3583
rect 2278 3538 2286 3569
rect 2215 3536 2286 3538
rect 2215 3535 2287 3536
rect 2098 3529 2109 3531
rect 2215 3530 2312 3535
rect 2278 3526 2312 3530
rect 2214 3502 2263 3510
rect 2192 3465 2200 3487
rect 2214 3493 2224 3502
rect 2255 3495 2263 3502
rect 2278 3494 2286 3526
rect 2301 3521 2312 3526
rect 2387 3523 2397 3556
rect 2301 3511 2342 3521
rect 2387 3514 2414 3523
rect 2387 3488 2397 3514
rect 2363 3461 2372 3477
rect 2363 3455 2398 3461
rect 1005 3422 1027 3428
rect 1054 3422 1867 3430
rect 1005 3416 1011 3422
rect 791 3399 832 3409
rect 877 3403 915 3411
rect 964 3410 1011 3416
rect 877 3402 914 3403
rect 877 3376 887 3402
rect 570 3347 605 3353
rect 853 3349 862 3365
rect 853 3343 888 3349
rect 903 3313 914 3402
rect 964 3398 971 3410
rect 1004 3398 1011 3410
rect 1054 3421 1858 3422
rect 1054 3398 1061 3421
rect 945 3378 951 3392
rect 985 3378 991 3392
rect 945 3373 1014 3378
rect 1036 3375 1042 3392
rect 608 3022 616 3027
rect 542 3016 616 3022
rect 542 3002 549 3016
rect 608 3000 616 3016
rect 748 3012 756 3020
rect 713 3006 756 3012
rect 564 2961 573 2992
rect 713 2992 721 3006
rect 627 2961 635 2992
rect 564 2959 635 2961
rect 564 2958 636 2959
rect 564 2953 661 2958
rect 627 2949 661 2953
rect 453 2917 460 2933
rect 563 2925 612 2933
rect 300 2888 309 2896
rect 470 2888 478 2908
rect 541 2891 549 2910
rect 563 2916 573 2925
rect 604 2918 612 2925
rect 627 2917 635 2949
rect 650 2944 661 2949
rect 736 2946 746 2979
rect 755 2946 1267 2947
rect 650 2934 691 2944
rect 736 2937 1267 2946
rect 736 2911 746 2937
rect 755 2936 1267 2937
rect 300 2881 462 2888
rect 300 2869 309 2881
rect 402 2880 440 2881
rect 298 2800 309 2869
rect 470 2877 617 2888
rect 712 2884 721 2900
rect 1259 2894 1267 2936
rect 1507 2923 1530 2929
rect 1507 2913 1513 2923
rect 1671 2913 1677 2929
rect 1259 2893 1523 2894
rect 1259 2887 1516 2893
rect 1522 2887 1523 2893
rect 1526 2891 1532 2904
rect 1547 2891 1553 2904
rect 1526 2885 1553 2891
rect 1567 2891 1573 2904
rect 1586 2891 1592 2904
rect 1567 2885 1592 2891
rect 1605 2891 1611 2904
rect 1629 2891 1635 2904
rect 1605 2885 1635 2891
rect 712 2878 747 2884
rect 1648 2882 1654 2904
rect 1689 2883 1696 2905
rect 1689 2882 1703 2883
rect 1776 2882 1844 2883
rect 470 2876 625 2877
rect 1648 2876 1662 2882
rect 1689 2877 1844 2882
rect 470 2866 478 2876
rect 1648 2870 1654 2876
rect 453 2847 460 2857
rect 608 2853 616 2858
rect 803 2857 811 2865
rect 542 2852 666 2853
rect 671 2852 679 2857
rect 542 2847 679 2852
rect 542 2833 549 2847
rect 608 2846 679 2847
rect 608 2831 616 2846
rect 671 2830 679 2846
rect 768 2851 811 2857
rect 1526 2864 1654 2870
rect 1526 2852 1533 2864
rect 768 2837 776 2851
rect 1566 2852 1573 2864
rect 1605 2853 1612 2864
rect 298 2773 308 2800
rect 564 2792 573 2823
rect 627 2792 635 2823
rect 564 2791 635 2792
rect 690 2791 698 2822
rect 564 2789 698 2791
rect 1507 2832 1513 2846
rect 1547 2832 1553 2846
rect 1647 2852 1654 2864
rect 1586 2832 1592 2845
rect 1689 2852 1696 2877
rect 1629 2832 1635 2845
rect 1507 2827 1635 2832
rect 1671 2829 1677 2846
rect 791 2791 801 2824
rect 806 2791 1557 2792
rect 564 2788 699 2789
rect 739 2788 746 2789
rect 564 2784 746 2788
rect 627 2780 746 2784
rect 690 2779 746 2780
rect 791 2782 1557 2791
rect 298 2770 309 2773
rect -1476 2396 -1450 2399
rect -1481 2395 55 2396
rect -1481 2394 69 2395
rect -1481 2370 42 2394
rect -1442 2369 -1352 2370
rect 14 2342 28 2356
rect -1389 2322 28 2342
rect -1421 2318 28 2322
rect -15 2249 -1 2286
rect -1335 2225 0 2249
rect -49 2195 -37 2212
rect -1307 2193 -37 2195
rect -1307 2184 -1298 2193
rect -1274 2184 -37 2193
rect -1307 2182 -37 2184
rect -120 2101 -91 2104
rect -1248 2099 -91 2101
rect -1220 2071 -91 2099
rect -541 2054 -136 2055
rect -1189 2053 -136 2054
rect -1167 2040 -136 2053
rect -1167 2039 -425 2040
rect -1136 1978 -181 1996
rect -281 1929 -252 1935
rect -1096 1905 -235 1929
rect -281 921 -252 1905
rect -281 -858 -252 903
rect -207 1321 -183 1978
rect -207 -790 -183 1307
rect -154 1745 -136 2040
rect -120 1994 -91 2071
rect -154 -513 -136 1728
rect -120 1607 -91 1973
rect -121 1593 -91 1607
rect -121 1147 -92 1593
rect -121 -42 -89 1147
rect -49 1106 -37 2182
rect -15 1586 -1 2225
rect -38 1097 -37 1106
rect -49 786 -37 1097
rect -49 -23 -36 786
rect -15 6 -1 1576
rect 14 1799 28 2318
rect 178 2232 202 2233
rect 14 37 28 1788
rect 167 2219 207 2232
rect 101 1728 111 1744
rect 86 1727 111 1728
rect 110 1307 132 1321
rect 147 1307 148 1321
rect 167 146 176 2219
rect 207 2094 215 2108
rect 275 1847 287 1848
rect 275 1800 287 1831
rect 196 1799 287 1800
rect 213 1788 287 1799
rect 196 1787 287 1788
rect 199 1576 248 1585
rect 249 1071 259 1514
rect 249 460 260 1071
rect 275 1019 287 1787
rect 300 1206 309 2770
rect 455 2755 462 2770
rect 563 2756 612 2764
rect 322 2719 464 2726
rect 472 2719 480 2746
rect 541 2723 549 2741
rect 563 2747 573 2756
rect 604 2749 612 2756
rect 627 2755 675 2763
rect 627 2748 635 2755
rect 667 2748 675 2755
rect 690 2747 698 2779
rect 791 2756 801 2782
rect 1839 2746 1844 2877
rect 2147 2814 2155 2818
rect 2147 2813 2265 2814
rect 2081 2809 2265 2813
rect 2081 2807 2155 2809
rect 2081 2793 2088 2807
rect 2147 2791 2155 2807
rect 2218 2808 2265 2809
rect 2218 2794 2225 2808
rect 2103 2752 2112 2783
rect 2166 2752 2174 2783
rect 2103 2750 2174 2752
rect 2281 2789 2288 2805
rect 2240 2753 2249 2784
rect 2298 2764 2306 2780
rect 2298 2763 2335 2764
rect 2298 2757 2317 2763
rect 2240 2750 2290 2753
rect 2103 2749 2175 2750
rect 2185 2749 2290 2750
rect 2103 2746 2290 2749
rect 767 2729 776 2745
rect 1839 2739 2092 2746
rect 2103 2745 2265 2746
rect 2103 2744 2249 2745
rect 2166 2743 2249 2744
rect 2166 2741 2187 2743
rect 767 2723 802 2729
rect 322 1498 330 2719
rect 402 2718 437 2719
rect 472 2708 617 2719
rect 2102 2716 2151 2724
rect 472 2707 625 2708
rect 472 2704 480 2707
rect 455 2685 462 2695
rect 588 2694 596 2699
rect 522 2693 646 2694
rect 651 2693 659 2698
rect 823 2696 831 2704
rect 522 2692 659 2693
rect 522 2691 714 2692
rect 719 2691 727 2696
rect 522 2688 727 2691
rect 522 2674 529 2688
rect 588 2687 727 2688
rect 588 2672 596 2687
rect 651 2685 727 2687
rect 651 2671 659 2685
rect 544 2633 553 2664
rect 719 2669 727 2685
rect 788 2690 831 2696
rect 788 2676 796 2690
rect 2080 2679 2088 2701
rect 2102 2707 2112 2716
rect 2143 2709 2151 2716
rect 2166 2718 2227 2727
rect 2252 2725 2260 2745
rect 2298 2738 2306 2757
rect 2166 2708 2174 2718
rect 2219 2709 2227 2718
rect 2239 2717 2265 2725
rect 2281 2719 2288 2729
rect 2239 2708 2249 2717
rect 607 2633 615 2664
rect 544 2632 615 2633
rect 670 2632 678 2663
rect 544 2630 678 2632
rect 738 2630 746 2661
rect 544 2629 679 2630
rect 694 2629 746 2630
rect 544 2628 746 2629
rect 811 2630 821 2663
rect 811 2629 1604 2630
rect 544 2627 747 2628
rect 759 2627 766 2628
rect 544 2625 766 2627
rect 607 2621 766 2625
rect 670 2620 766 2621
rect 702 2619 766 2620
rect 738 2618 766 2619
rect 811 2622 1595 2629
rect 1602 2622 1604 2629
rect 811 2621 838 2622
rect 454 2600 461 2616
rect 543 2597 592 2605
rect 400 2571 435 2572
rect 341 2564 463 2571
rect 471 2569 479 2591
rect 341 1817 349 2564
rect 471 2560 503 2569
rect 521 2564 529 2582
rect 543 2588 553 2597
rect 584 2590 592 2597
rect 607 2596 655 2604
rect 670 2602 678 2603
rect 607 2589 615 2596
rect 647 2589 655 2596
rect 669 2595 723 2602
rect 670 2588 678 2595
rect 702 2594 723 2595
rect 715 2587 723 2594
rect 738 2586 746 2618
rect 811 2595 821 2621
rect 787 2568 796 2584
rect 787 2562 822 2568
rect 471 2559 597 2560
rect 471 2549 479 2559
rect 495 2549 597 2559
rect 1141 2557 1281 2558
rect 1141 2555 1265 2557
rect 496 2548 605 2549
rect 763 2546 1265 2555
rect 1280 2546 1281 2557
rect 763 2545 1281 2546
rect 454 2530 461 2540
rect 2869 2537 2878 3601
rect 2928 2606 2937 4189
rect 2972 2915 2982 5628
rect 3023 5624 3028 5665
rect 3050 5668 3080 5674
rect 3103 5668 3166 5674
rect 3050 5653 3058 5668
rect 3033 5634 3040 5644
rect 3107 5624 3115 5668
rect 3023 5617 3125 5624
rect 3158 3183 3165 5668
rect 3204 5646 3218 5677
rect 2972 2902 2982 2903
rect 2928 2582 2937 2592
rect 2869 2513 2878 2523
rect 793 2504 1293 2506
rect 793 2494 795 2504
rect 804 2494 1293 2504
rect 793 2493 1308 2494
rect 597 2475 605 2480
rect 531 2474 655 2475
rect 660 2474 668 2479
rect 531 2473 668 2474
rect 531 2472 723 2473
rect 728 2472 736 2477
rect 893 2476 901 2484
rect 787 2472 795 2476
rect 531 2469 795 2472
rect 531 2455 538 2469
rect 597 2468 795 2469
rect 597 2453 605 2468
rect 660 2466 795 2468
rect 660 2452 668 2466
rect 726 2465 795 2466
rect 388 2411 400 2422
rect 553 2414 562 2445
rect 728 2450 736 2465
rect 616 2414 624 2445
rect 553 2413 624 2414
rect 679 2413 687 2444
rect 787 2449 795 2465
rect 858 2470 901 2476
rect 858 2456 866 2470
rect 553 2411 687 2413
rect 747 2411 755 2442
rect 553 2410 688 2411
rect 703 2410 755 2411
rect 806 2410 814 2441
rect 553 2408 814 2410
rect 881 2410 891 2443
rect 895 2410 1639 2412
rect 553 2407 815 2408
rect 827 2407 836 2408
rect 553 2406 836 2407
rect 616 2402 836 2406
rect 679 2401 836 2402
rect 711 2400 836 2401
rect 747 2399 836 2400
rect 806 2398 836 2399
rect 881 2402 1639 2410
rect 881 2401 908 2402
rect 1645 2402 1698 2412
rect 454 2368 461 2384
rect 552 2378 601 2386
rect 471 2342 479 2359
rect 504 2342 512 2343
rect 530 2342 538 2363
rect 552 2369 562 2378
rect 593 2371 601 2378
rect 616 2377 664 2385
rect 679 2383 687 2384
rect 616 2370 624 2377
rect 656 2370 664 2377
rect 678 2376 732 2383
rect 679 2369 687 2376
rect 711 2375 732 2376
rect 724 2368 732 2375
rect 747 2381 755 2382
rect 770 2381 791 2382
rect 747 2374 791 2381
rect 747 2367 755 2374
rect 783 2367 791 2374
rect 806 2366 814 2398
rect 881 2375 891 2401
rect 857 2348 866 2364
rect 857 2342 892 2348
rect 471 2341 556 2342
rect 395 2339 437 2340
rect 370 2332 463 2339
rect 372 2232 382 2332
rect 471 2331 606 2341
rect 471 2317 479 2331
rect 504 2330 606 2331
rect 1067 2338 1279 2339
rect 1067 2337 1263 2338
rect 852 2336 1263 2337
rect 505 2329 614 2330
rect 772 2326 1263 2336
rect 454 2298 461 2308
rect 381 2219 382 2232
rect 372 2116 382 2219
rect 372 2104 382 2108
rect 742 2107 1001 2109
rect 428 2096 727 2106
rect 742 2100 993 2107
rect 1000 2100 1001 2107
rect 742 2099 1001 2100
rect 477 2085 485 2096
rect 680 2085 688 2096
rect 411 2079 485 2085
rect 411 2065 418 2079
rect 477 2063 485 2079
rect 614 2079 688 2085
rect 614 2065 621 2079
rect 433 2024 442 2055
rect 680 2063 688 2079
rect 496 2034 504 2055
rect 495 2024 504 2034
rect 433 2021 504 2024
rect 636 2024 645 2055
rect 699 2024 707 2055
rect 636 2023 707 2024
rect 743 2023 752 2099
rect 867 2085 875 2094
rect 1048 2085 1056 2094
rect 801 2079 875 2085
rect 801 2065 808 2079
rect 867 2063 875 2079
rect 433 2016 530 2021
rect 636 2016 752 2023
rect 982 2079 1056 2085
rect 982 2065 989 2079
rect 823 2024 832 2055
rect 1048 2063 1056 2079
rect 886 2024 894 2055
rect 823 2023 894 2024
rect 1004 2024 1013 2055
rect 1067 2024 1075 2055
rect 1139 2050 1146 2066
rect 1156 2025 1164 2041
rect 1004 2023 1075 2024
rect 1081 2023 1148 2025
rect 823 2016 940 2023
rect 1004 2016 1148 2023
rect 1156 2016 1507 2025
rect 496 2012 530 2016
rect 432 1988 481 1996
rect 410 1951 418 1973
rect 432 1979 442 1988
rect 473 1981 481 1988
rect 496 1980 504 2012
rect 519 1939 530 2012
rect 699 2014 752 2016
rect 886 2014 940 2016
rect 635 1988 684 1996
rect 613 1951 621 1973
rect 635 1979 645 1988
rect 676 1981 684 1988
rect 699 1980 707 2014
rect 822 1988 871 1996
rect 800 1951 808 1973
rect 822 1979 832 1988
rect 863 1981 871 1988
rect 886 1980 894 2014
rect 519 1938 876 1939
rect 519 1930 689 1938
rect 696 1931 876 1938
rect 883 1931 917 1939
rect 696 1930 917 1931
rect 519 1928 917 1930
rect 928 1920 940 2014
rect 1067 2014 1095 2016
rect 1003 1988 1052 1996
rect 981 1951 989 1973
rect 1003 1979 1013 1988
rect 1044 1981 1052 1988
rect 1067 1980 1075 2014
rect 1156 1999 1164 2016
rect 1139 1980 1146 1990
rect 928 1913 1057 1920
rect 1064 1913 1097 1920
rect 928 1910 1097 1913
rect 748 1818 1007 1820
rect 351 1804 361 1815
rect 434 1807 733 1817
rect 748 1811 999 1818
rect 1006 1811 1007 1818
rect 748 1810 1007 1811
rect 483 1796 491 1807
rect 686 1796 694 1807
rect 417 1790 491 1796
rect 417 1776 424 1790
rect 483 1774 491 1790
rect 620 1790 694 1796
rect 620 1776 627 1790
rect 439 1735 448 1766
rect 686 1774 694 1790
rect 502 1745 510 1766
rect 501 1735 510 1745
rect 439 1732 510 1735
rect 642 1735 651 1766
rect 705 1735 713 1766
rect 642 1734 713 1735
rect 749 1734 758 1810
rect 873 1796 881 1805
rect 1054 1796 1062 1805
rect 807 1790 881 1796
rect 807 1776 814 1790
rect 873 1774 881 1790
rect 439 1727 536 1732
rect 642 1727 758 1734
rect 988 1790 1062 1796
rect 988 1776 995 1790
rect 829 1735 838 1766
rect 1054 1774 1062 1790
rect 892 1735 900 1766
rect 829 1734 900 1735
rect 1010 1735 1019 1766
rect 1073 1735 1081 1766
rect 1141 1758 1148 1774
rect 1010 1734 1081 1735
rect 1099 1734 1128 1735
rect 829 1727 946 1734
rect 1010 1733 1128 1734
rect 1158 1733 1166 1749
rect 1010 1727 1150 1733
rect 502 1723 536 1727
rect 438 1699 487 1707
rect 416 1662 424 1684
rect 438 1690 448 1699
rect 479 1692 487 1699
rect 502 1691 510 1723
rect 525 1650 536 1723
rect 705 1725 758 1727
rect 892 1725 946 1727
rect 641 1699 690 1707
rect 619 1662 627 1684
rect 641 1690 651 1699
rect 682 1692 690 1699
rect 705 1691 713 1725
rect 828 1699 877 1707
rect 806 1662 814 1684
rect 828 1690 838 1699
rect 869 1692 877 1699
rect 892 1691 900 1725
rect 525 1649 882 1650
rect 525 1641 695 1649
rect 702 1642 882 1649
rect 889 1642 923 1650
rect 702 1641 923 1642
rect 525 1639 923 1641
rect 934 1631 946 1725
rect 1073 1725 1150 1727
rect 1009 1699 1058 1707
rect 987 1662 995 1684
rect 1009 1690 1019 1699
rect 1050 1692 1058 1699
rect 1073 1691 1081 1725
rect 1099 1724 1150 1725
rect 1158 1724 1191 1733
rect 1158 1707 1166 1724
rect 1141 1688 1148 1698
rect 1178 1649 1189 1724
rect 934 1624 1063 1631
rect 1070 1624 1103 1631
rect 934 1621 1103 1624
rect 1179 1510 1188 1649
rect 1426 1512 1434 1516
rect 1563 1512 1571 1517
rect 2147 1515 2155 1519
rect 2147 1514 2265 1515
rect 1426 1511 1571 1512
rect 768 1501 1027 1503
rect 1179 1502 1294 1510
rect 1307 1502 1309 1510
rect 322 1496 380 1498
rect 328 1489 380 1496
rect 322 1488 380 1489
rect 454 1490 753 1500
rect 768 1494 1019 1501
rect 1026 1494 1027 1501
rect 768 1493 1027 1494
rect 503 1479 511 1490
rect 706 1479 714 1490
rect 437 1473 511 1479
rect 437 1459 444 1473
rect 503 1457 511 1473
rect 640 1473 714 1479
rect 640 1459 647 1473
rect 459 1418 468 1449
rect 706 1457 714 1473
rect 522 1428 530 1449
rect 521 1418 530 1428
rect 459 1415 530 1418
rect 662 1418 671 1449
rect 725 1418 733 1449
rect 662 1417 733 1418
rect 769 1417 778 1493
rect 893 1479 901 1488
rect 1074 1479 1082 1488
rect 827 1473 901 1479
rect 827 1459 834 1473
rect 893 1457 901 1473
rect 459 1410 556 1415
rect 662 1410 778 1417
rect 1008 1473 1082 1479
rect 1008 1459 1015 1473
rect 849 1418 858 1449
rect 1074 1457 1082 1473
rect 912 1418 920 1449
rect 849 1417 920 1418
rect 1030 1418 1039 1449
rect 1093 1418 1101 1449
rect 1166 1441 1173 1457
rect 1302 1437 1309 1502
rect 1360 1507 1571 1511
rect 1360 1505 1434 1507
rect 1360 1491 1367 1505
rect 1426 1489 1434 1505
rect 1497 1506 1571 1507
rect 1497 1492 1504 1506
rect 1382 1450 1391 1481
rect 1563 1490 1571 1506
rect 2081 1510 2265 1514
rect 2081 1508 2155 1510
rect 2081 1494 2088 1508
rect 1445 1450 1453 1481
rect 1382 1448 1453 1450
rect 1519 1451 1528 1482
rect 1582 1451 1590 1482
rect 1628 1477 1635 1493
rect 2147 1492 2155 1508
rect 2218 1509 2265 1510
rect 2218 1495 2225 1509
rect 1519 1449 1590 1451
rect 1645 1450 1653 1468
rect 2103 1453 2112 1484
rect 2166 1453 2174 1484
rect 2103 1451 2174 1453
rect 2281 1490 2288 1506
rect 2240 1454 2249 1485
rect 2298 1458 2306 1481
rect 2298 1454 3088 1458
rect 2240 1451 2290 1454
rect 2103 1450 2175 1451
rect 2185 1450 2290 1451
rect 1519 1448 1591 1449
rect 1645 1448 1841 1450
rect 1382 1447 1454 1448
rect 1464 1447 1637 1448
rect 1382 1443 1637 1447
rect 1382 1442 1528 1443
rect 1445 1441 1528 1442
rect 1445 1439 1466 1441
rect 1582 1439 1637 1443
rect 1030 1417 1101 1418
rect 849 1410 966 1417
rect 1030 1416 1136 1417
rect 1183 1416 1191 1432
rect 1302 1428 1371 1437
rect 1377 1428 1380 1437
rect 1235 1416 1309 1417
rect 1030 1410 1175 1416
rect 522 1406 556 1410
rect 458 1382 507 1390
rect 436 1345 444 1367
rect 458 1373 468 1382
rect 499 1375 507 1382
rect 522 1374 530 1406
rect 545 1333 556 1406
rect 725 1408 778 1410
rect 912 1408 966 1410
rect 661 1382 710 1390
rect 639 1345 647 1367
rect 661 1373 671 1382
rect 702 1375 710 1382
rect 725 1374 733 1408
rect 848 1382 897 1390
rect 826 1345 834 1367
rect 848 1373 858 1382
rect 889 1375 897 1382
rect 912 1374 920 1408
rect 545 1332 902 1333
rect 545 1324 715 1332
rect 722 1325 902 1332
rect 909 1325 943 1333
rect 722 1324 943 1325
rect 545 1322 943 1324
rect 954 1314 966 1408
rect 1093 1408 1175 1410
rect 1029 1382 1078 1390
rect 1007 1345 1015 1367
rect 1029 1373 1039 1382
rect 1070 1375 1078 1382
rect 1093 1374 1101 1408
rect 1110 1407 1175 1408
rect 1183 1407 1263 1416
rect 1277 1407 1309 1416
rect 1183 1390 1191 1407
rect 1166 1371 1173 1381
rect 1302 1339 1309 1407
rect 1381 1414 1430 1422
rect 1359 1377 1367 1399
rect 1381 1405 1391 1414
rect 1422 1407 1430 1414
rect 1445 1416 1506 1425
rect 1445 1406 1453 1416
rect 1498 1407 1506 1416
rect 1518 1415 1567 1423
rect 1518 1406 1528 1415
rect 1559 1408 1567 1415
rect 1582 1407 1590 1439
rect 1598 1438 1637 1439
rect 1645 1447 1969 1448
rect 2103 1447 2290 1450
rect 1645 1440 2092 1447
rect 2103 1446 2265 1447
rect 2103 1445 2259 1446
rect 2166 1444 2259 1445
rect 2166 1442 2187 1444
rect 1645 1426 1653 1440
rect 1829 1439 1969 1440
rect 2102 1417 2151 1425
rect 1628 1407 1635 1417
rect 2080 1380 2088 1402
rect 2102 1408 2112 1417
rect 2143 1410 2151 1417
rect 2166 1419 2227 1428
rect 2251 1426 2259 1444
rect 2298 1439 2306 1454
rect 2166 1409 2174 1419
rect 2219 1410 2227 1419
rect 2239 1418 2265 1426
rect 2281 1420 2288 1430
rect 2239 1409 2249 1418
rect 1302 1328 1572 1339
rect 1579 1328 1582 1339
rect 954 1307 1083 1314
rect 1090 1307 1123 1314
rect 954 1304 1123 1307
rect 766 1210 1025 1212
rect 300 1196 382 1206
rect 452 1199 751 1209
rect 766 1203 1017 1210
rect 1024 1203 1025 1210
rect 766 1202 1025 1203
rect 285 1001 287 1019
rect 358 976 368 1196
rect 501 1188 509 1199
rect 704 1188 712 1199
rect 435 1182 509 1188
rect 435 1168 442 1182
rect 501 1166 509 1182
rect 638 1182 712 1188
rect 638 1168 645 1182
rect 457 1127 466 1158
rect 704 1166 712 1182
rect 520 1137 528 1158
rect 519 1127 528 1137
rect 457 1124 528 1127
rect 660 1127 669 1158
rect 723 1127 731 1158
rect 660 1126 731 1127
rect 767 1126 776 1202
rect 891 1188 899 1197
rect 1072 1188 1080 1197
rect 825 1182 899 1188
rect 825 1168 832 1182
rect 891 1166 899 1182
rect 457 1119 554 1124
rect 660 1119 776 1126
rect 1006 1182 1080 1188
rect 1006 1168 1013 1182
rect 847 1127 856 1158
rect 1072 1166 1080 1182
rect 910 1127 918 1158
rect 847 1126 918 1127
rect 1028 1127 1037 1158
rect 1091 1127 1099 1158
rect 1175 1150 1182 1166
rect 1028 1126 1099 1127
rect 847 1119 964 1126
rect 1028 1125 1119 1126
rect 1192 1125 1200 1141
rect 1235 1125 1252 1126
rect 1028 1119 1184 1125
rect 520 1115 554 1119
rect 456 1091 505 1099
rect 434 1054 442 1076
rect 456 1082 466 1091
rect 497 1084 505 1091
rect 520 1083 528 1115
rect 543 1042 554 1115
rect 723 1117 776 1119
rect 910 1117 964 1119
rect 659 1091 708 1099
rect 637 1054 645 1076
rect 659 1082 669 1091
rect 700 1084 708 1091
rect 723 1083 731 1117
rect 846 1091 895 1099
rect 824 1054 832 1076
rect 846 1082 856 1091
rect 887 1084 895 1091
rect 910 1083 918 1117
rect 543 1041 900 1042
rect 543 1033 713 1041
rect 720 1034 900 1041
rect 907 1034 941 1042
rect 720 1033 941 1034
rect 543 1031 941 1033
rect 952 1023 964 1117
rect 1091 1117 1184 1119
rect 1027 1091 1076 1099
rect 1005 1054 1013 1076
rect 1027 1082 1037 1091
rect 1068 1084 1076 1091
rect 1091 1083 1099 1117
rect 1153 1116 1184 1117
rect 1192 1116 1236 1125
rect 1250 1124 1443 1125
rect 1250 1117 1435 1124
rect 1250 1116 1252 1117
rect 1192 1099 1200 1116
rect 1175 1080 1182 1090
rect 952 1016 1081 1023
rect 1088 1016 1121 1023
rect 952 1013 1121 1016
rect 358 692 368 962
rect 554 756 562 761
rect 488 750 562 756
rect 488 736 495 750
rect 554 734 562 750
rect 694 746 702 754
rect 659 740 702 746
rect 510 695 519 726
rect 659 726 667 740
rect 573 695 581 726
rect 510 693 581 695
rect 510 692 582 693
rect 357 691 410 692
rect 357 679 383 691
rect 409 679 410 691
rect 510 687 607 692
rect 357 677 410 679
rect 573 683 607 687
rect 399 651 406 667
rect 509 659 558 667
rect 416 622 424 642
rect 487 625 495 644
rect 509 650 519 659
rect 550 652 558 659
rect 573 651 581 683
rect 596 678 607 683
rect 682 680 692 713
rect 2147 684 2155 688
rect 2147 683 2265 684
rect 701 680 1268 681
rect 596 668 637 678
rect 682 671 1268 680
rect 682 645 692 671
rect 701 670 1268 671
rect 977 669 1035 670
rect 392 615 408 622
rect 383 614 386 615
rect 416 611 563 622
rect 658 618 667 634
rect 1260 628 1268 670
rect 2081 679 2265 683
rect 2081 677 2155 679
rect 2081 663 2088 677
rect 1567 657 1590 663
rect 1567 647 1573 657
rect 1731 647 1737 663
rect 2147 661 2155 677
rect 1260 627 1583 628
rect 1260 621 1576 627
rect 1582 621 1583 627
rect 1586 625 1592 638
rect 1607 625 1613 638
rect 1586 619 1613 625
rect 1627 625 1633 638
rect 1646 625 1652 638
rect 1627 619 1652 625
rect 1665 625 1671 638
rect 1689 625 1695 638
rect 1665 619 1695 625
rect 2218 678 2265 679
rect 2218 664 2225 678
rect 658 612 693 618
rect 1708 616 1714 638
rect 1749 617 1756 639
rect 2103 622 2112 653
rect 2166 622 2174 653
rect 2103 620 2174 622
rect 2281 659 2288 675
rect 2240 623 2249 654
rect 2298 626 2306 650
rect 2240 620 2290 623
rect 2103 619 2175 620
rect 2185 619 2290 620
rect 1749 616 1763 617
rect 1836 616 2051 617
rect 2103 616 2290 619
rect 2298 619 3063 626
rect 416 610 571 611
rect 1708 610 1722 616
rect 1749 611 2092 616
rect 416 600 424 610
rect 1708 604 1714 610
rect 399 581 406 591
rect 554 587 562 592
rect 749 591 757 599
rect 488 586 612 587
rect 617 586 625 591
rect 488 581 625 586
rect 488 567 495 581
rect 554 580 625 581
rect 554 565 562 580
rect 617 564 625 580
rect 714 585 757 591
rect 1586 598 1714 604
rect 1586 586 1593 598
rect 714 571 722 585
rect 1626 586 1633 598
rect 1665 587 1672 598
rect 510 526 519 557
rect 573 526 581 557
rect 510 525 581 526
rect 636 525 644 556
rect 510 523 644 525
rect 1567 566 1573 580
rect 1607 566 1613 580
rect 1707 586 1714 598
rect 1646 566 1652 579
rect 1749 586 1756 611
rect 2036 609 2092 611
rect 2103 615 2265 616
rect 2103 614 2249 615
rect 2166 613 2249 614
rect 2166 611 2187 613
rect 2102 586 2151 594
rect 1689 566 1695 579
rect 1567 561 1695 566
rect 1731 563 1737 580
rect 737 525 747 558
rect 2080 549 2088 571
rect 2102 577 2112 586
rect 2143 579 2151 586
rect 2166 588 2227 597
rect 2252 595 2260 615
rect 2298 608 2306 619
rect 2166 578 2174 588
rect 2219 579 2227 588
rect 2239 587 2265 595
rect 2281 589 2288 599
rect 2239 578 2249 587
rect 752 525 1325 526
rect 1496 525 1617 526
rect 286 521 364 523
rect 303 512 364 521
rect 286 510 364 512
rect 510 522 645 523
rect 685 522 692 523
rect 510 518 692 522
rect 573 514 692 518
rect 636 513 692 514
rect 737 517 1617 525
rect 737 516 1325 517
rect 1496 516 1617 517
rect 401 489 408 504
rect 509 490 558 498
rect 249 453 410 460
rect 418 453 426 480
rect 487 457 495 475
rect 509 481 519 490
rect 550 483 558 490
rect 573 489 621 497
rect 573 482 581 489
rect 613 482 621 489
rect 636 481 644 513
rect 737 490 747 516
rect 713 463 722 479
rect 713 457 748 463
rect 418 442 563 453
rect 418 441 571 442
rect 418 438 426 441
rect 401 419 408 429
rect 534 428 542 433
rect 468 427 592 428
rect 597 427 605 432
rect 769 430 777 438
rect 468 426 605 427
rect 468 425 660 426
rect 665 425 673 430
rect 468 422 673 425
rect 468 408 475 422
rect 534 421 673 422
rect 534 406 542 421
rect 597 419 673 421
rect 597 405 605 419
rect 351 367 383 368
rect 490 367 499 398
rect 665 403 673 419
rect 734 424 777 430
rect 734 410 742 424
rect 553 367 561 398
rect 351 351 364 367
rect 490 366 561 367
rect 616 366 624 397
rect 490 364 624 366
rect 684 364 692 395
rect 490 363 625 364
rect 640 363 692 364
rect 490 362 692 363
rect 757 364 767 397
rect 757 363 1325 364
rect 1496 363 1664 364
rect 490 361 693 362
rect 705 361 712 362
rect 490 359 712 361
rect 553 355 712 359
rect 616 354 712 355
rect 648 353 712 354
rect 684 352 712 353
rect 757 356 1655 363
rect 1662 356 1664 363
rect 757 355 784 356
rect 1306 355 1566 356
rect 400 334 407 350
rect 489 331 538 339
rect 378 305 381 306
rect 378 299 409 305
rect 364 298 409 299
rect 417 303 425 325
rect 417 294 449 303
rect 467 298 475 316
rect 489 322 499 331
rect 530 324 538 331
rect 553 330 601 338
rect 616 336 624 337
rect 553 323 561 330
rect 593 323 601 330
rect 615 329 669 336
rect 616 322 624 329
rect 648 328 669 329
rect 661 321 669 328
rect 684 320 692 352
rect 757 329 767 355
rect 733 302 742 318
rect 733 296 768 302
rect 417 293 543 294
rect 417 283 425 293
rect 441 283 543 293
rect 1142 291 1282 292
rect 1142 289 1266 291
rect 442 282 551 283
rect 709 280 1266 289
rect 1281 280 1282 291
rect 709 279 1282 280
rect 400 264 407 274
rect 739 238 1294 240
rect 739 228 741 238
rect 750 228 1294 238
rect 739 227 1309 228
rect 543 209 551 214
rect 477 208 601 209
rect 606 208 614 213
rect 477 207 614 208
rect 477 206 669 207
rect 674 206 682 211
rect 839 210 847 218
rect 733 206 741 210
rect 477 203 741 206
rect 477 189 484 203
rect 543 202 741 203
rect 543 187 551 202
rect 606 200 741 202
rect 606 186 614 200
rect 672 199 741 200
rect 499 148 508 179
rect 674 184 682 199
rect 562 148 570 179
rect 499 147 570 148
rect 625 147 633 178
rect 733 183 741 199
rect 804 204 847 210
rect 804 190 812 204
rect 167 145 377 146
rect 499 145 633 147
rect 693 145 701 176
rect 167 132 364 145
rect 499 144 634 145
rect 649 144 701 145
rect 752 144 760 175
rect 499 142 760 144
rect 827 144 837 177
rect 841 144 1325 146
rect 1496 144 1699 146
rect 499 141 761 142
rect 773 141 782 142
rect 499 140 782 141
rect 562 136 782 140
rect 625 135 782 136
rect 657 134 782 135
rect 693 133 782 134
rect 752 132 782 133
rect 827 136 1699 144
rect 827 135 854 136
rect 167 131 377 132
rect 400 102 407 118
rect 498 112 547 120
rect 417 76 425 93
rect 450 76 458 77
rect 476 76 484 97
rect 498 103 508 112
rect 539 105 547 112
rect 562 111 610 119
rect 625 117 633 118
rect 562 104 570 111
rect 602 104 610 111
rect 624 110 678 117
rect 625 103 633 110
rect 657 109 678 110
rect 670 102 678 109
rect 693 115 701 116
rect 716 115 737 116
rect 693 108 737 115
rect 693 101 701 108
rect 729 101 737 108
rect 752 100 760 132
rect 827 109 837 135
rect 1001 134 1048 136
rect 1705 136 1758 146
rect 803 82 812 98
rect 803 76 838 82
rect 231 74 255 75
rect 68 73 383 74
rect 68 67 409 73
rect 45 66 409 67
rect 417 72 470 76
rect 491 75 502 76
rect 491 72 552 75
rect 14 34 136 37
rect 14 23 137 34
rect -15 -11 93 6
rect -15 -12 -1 -11
rect 44 -23 57 -22
rect -50 -34 57 -23
rect -118 -458 -89 -42
rect -118 -486 -89 -472
rect -137 -527 -136 -513
rect -207 -814 -183 -805
rect 44 -825 57 -34
rect 78 -759 92 -11
rect 118 -484 137 23
rect 231 -431 255 66
rect 417 65 552 72
rect 417 51 425 65
rect 450 64 552 65
rect 1013 72 1280 73
rect 1013 71 1264 72
rect 798 70 1264 71
rect 718 60 1264 70
rect 400 32 407 42
rect 3203 -255 3218 5646
rect 3277 5594 3288 5677
rect 3304 5627 3311 5643
rect 3277 5588 3278 5594
rect 3321 5597 3329 5618
rect 3358 5597 3368 5598
rect 3321 5591 3368 5597
rect 3321 5576 3329 5591
rect 3304 5557 3311 5567
rect 3356 5534 3367 5591
rect 3236 3690 5321 3699
rect 5328 3690 5661 3699
rect 4453 2606 4896 2607
rect 4462 2604 4896 2606
rect 4462 2592 4881 2604
rect 4435 2590 4881 2592
rect 4888 2590 4896 2604
rect 4495 2523 5138 2537
rect 5145 2523 5149 2537
rect 4477 2522 5098 2523
rect 3407 1454 4858 1458
rect 4840 1032 4846 1454
rect 5047 1043 5070 1049
rect 5047 1033 5053 1043
rect 5170 1033 5176 1049
rect 4790 1006 4813 1012
rect 4790 996 4796 1006
rect 4913 996 4919 1012
rect 5066 1011 5072 1024
rect 5087 1011 5093 1024
rect 5066 1005 5093 1011
rect 5104 1011 5110 1024
rect 5128 1011 5134 1024
rect 5104 1005 5134 1011
rect 4809 974 4815 987
rect 4830 974 4836 987
rect 4809 968 4836 974
rect 4847 974 4853 987
rect 4871 974 4877 987
rect 4847 968 4877 974
rect 5147 1002 5153 1024
rect 5188 1003 5195 1025
rect 5147 996 5161 1002
rect 5188 997 5202 1003
rect 4890 965 4896 987
rect 5147 990 5153 996
rect 4931 966 4938 988
rect 5066 984 5153 990
rect 5066 972 5073 984
rect 5104 973 5111 984
rect 5146 972 5153 984
rect 4890 959 4904 965
rect 4931 960 4945 966
rect 4890 953 4896 959
rect 4809 947 4896 953
rect 4809 935 4816 947
rect 4847 936 4854 947
rect 4889 935 4896 947
rect 4790 915 4796 929
rect 4830 915 4836 929
rect 4931 935 4938 960
rect 5047 952 5053 966
rect 5087 952 5093 966
rect 5188 972 5195 997
rect 5128 952 5134 965
rect 5047 947 5134 952
rect 5170 949 5176 966
rect 4871 915 4877 928
rect 4790 910 4877 915
rect 4913 912 4919 929
rect 4546 851 4569 857
rect 4546 841 4552 851
rect 4669 841 4675 857
rect 4565 819 4571 832
rect 4586 819 4592 832
rect 4565 813 4592 819
rect 4603 819 4609 832
rect 4627 819 4633 832
rect 4603 813 4633 819
rect 4646 810 4652 832
rect 4687 811 4694 833
rect 4646 804 4660 810
rect 4687 805 4701 811
rect 4646 798 4652 804
rect 4565 792 4652 798
rect 4565 780 4572 792
rect 4603 781 4610 792
rect 4645 780 4652 792
rect 4546 760 4552 774
rect 4586 760 4592 774
rect 4687 780 4694 805
rect 4627 760 4633 773
rect 4546 755 4633 760
rect 4669 757 4675 774
rect 5248 670 5271 676
rect 5248 660 5254 670
rect 5339 660 5345 676
rect 5267 638 5273 651
rect 5288 638 5294 651
rect 5267 632 5294 638
rect 5308 629 5314 651
rect 5357 630 5364 652
rect 3834 619 5095 626
rect 3827 618 5095 619
rect 5104 618 5110 626
rect 5308 623 5330 629
rect 5357 624 5371 630
rect 5308 617 5314 623
rect 5267 611 5314 617
rect 5267 599 5274 611
rect 5307 599 5314 611
rect 5357 599 5364 624
rect 5248 579 5254 593
rect 5288 579 5294 593
rect 5248 574 5317 579
rect 5339 576 5345 593
rect 3203 -272 3218 -267
rect 760 -291 768 -286
rect 694 -297 768 -291
rect 694 -311 701 -297
rect 760 -313 768 -297
rect 900 -301 908 -293
rect 865 -307 908 -301
rect 716 -352 725 -321
rect 865 -321 873 -307
rect 779 -352 787 -321
rect 716 -354 787 -352
rect 1348 -333 1356 -329
rect 1348 -334 1466 -333
rect 716 -355 788 -354
rect 716 -360 813 -355
rect 779 -364 813 -360
rect 715 -388 764 -380
rect 693 -425 701 -403
rect 715 -397 725 -388
rect 756 -395 764 -388
rect 779 -396 787 -364
rect 802 -369 813 -364
rect 888 -367 898 -334
rect 1282 -338 1466 -334
rect 1282 -340 1356 -338
rect 1282 -354 1289 -340
rect 1348 -356 1356 -340
rect 1419 -339 1466 -338
rect 1419 -353 1426 -339
rect 802 -379 843 -369
rect 888 -376 1187 -367
rect 888 -402 898 -376
rect 909 -377 1187 -376
rect 1179 -400 1187 -377
rect 1304 -395 1313 -364
rect 1367 -395 1375 -364
rect 1304 -397 1375 -395
rect 1482 -358 1489 -342
rect 1441 -394 1450 -363
rect 1441 -397 1491 -394
rect 1304 -398 1376 -397
rect 1386 -398 1491 -397
rect 1179 -401 1267 -400
rect 1304 -401 1491 -398
rect 1499 -395 1507 -367
rect 1499 -399 4555 -395
rect 1179 -408 1293 -401
rect 1304 -402 1466 -401
rect 1304 -403 1450 -402
rect 1367 -404 1450 -403
rect 1367 -406 1388 -404
rect 1179 -409 1267 -408
rect 1179 -411 1187 -409
rect 864 -429 873 -413
rect 200 -432 352 -431
rect 200 -445 335 -432
rect 864 -435 899 -429
rect 1303 -431 1352 -423
rect 217 -472 397 -458
rect 330 -473 397 -472
rect 413 -473 414 -458
rect 467 -475 468 -466
rect 1281 -468 1289 -446
rect 1303 -440 1313 -431
rect 1344 -438 1352 -431
rect 1367 -429 1428 -420
rect 1454 -422 1462 -402
rect 1499 -409 1507 -399
rect 1367 -439 1375 -429
rect 1420 -438 1428 -429
rect 1440 -430 1466 -422
rect 1482 -428 1489 -418
rect 1440 -439 1450 -430
rect 467 -483 481 -475
rect 327 -484 482 -483
rect 118 -498 482 -484
rect 762 -489 770 -484
rect 696 -495 770 -489
rect 696 -509 703 -495
rect 219 -527 485 -514
rect 762 -511 770 -495
rect 902 -499 910 -491
rect 219 -528 352 -527
rect 471 -636 485 -527
rect 867 -505 910 -499
rect 718 -550 727 -519
rect 867 -519 875 -505
rect 781 -550 789 -519
rect 718 -552 789 -550
rect 1348 -523 1356 -519
rect 1348 -524 1466 -523
rect 718 -553 790 -552
rect 718 -558 815 -553
rect 781 -562 815 -558
rect 717 -586 766 -578
rect 695 -623 703 -601
rect 717 -595 727 -586
rect 758 -593 766 -586
rect 781 -594 789 -562
rect 804 -567 815 -562
rect 890 -565 900 -532
rect 1282 -528 1466 -524
rect 1282 -530 1356 -528
rect 1282 -544 1289 -530
rect 1348 -546 1356 -530
rect 1419 -529 1466 -528
rect 1419 -543 1426 -529
rect 972 -557 980 -555
rect 972 -565 1187 -557
rect 890 -567 1187 -565
rect 804 -577 845 -567
rect 890 -574 981 -567
rect 890 -600 900 -574
rect 1179 -590 1187 -567
rect 1304 -585 1313 -554
rect 1367 -585 1375 -554
rect 1304 -587 1375 -585
rect 1482 -548 1489 -532
rect 1441 -584 1450 -553
rect 1441 -587 1491 -584
rect 1304 -588 1376 -587
rect 1386 -588 1491 -587
rect 1179 -591 1267 -590
rect 1304 -591 1491 -588
rect 1499 -586 1507 -557
rect 1499 -590 4799 -586
rect 1179 -598 1293 -591
rect 1304 -592 1466 -591
rect 1304 -593 1450 -592
rect 1367 -594 1450 -593
rect 1367 -596 1388 -594
rect 1179 -599 1267 -598
rect 1179 -601 1187 -599
rect 866 -627 875 -611
rect 1303 -621 1352 -613
rect 866 -633 901 -627
rect 471 -646 485 -645
rect 1281 -658 1289 -636
rect 1303 -630 1313 -621
rect 1344 -628 1352 -621
rect 1367 -619 1428 -610
rect 1455 -612 1463 -592
rect 1499 -599 1507 -590
rect 1367 -629 1375 -619
rect 1420 -628 1428 -619
rect 1440 -620 1466 -612
rect 1482 -618 1489 -608
rect 1440 -629 1450 -620
rect 762 -687 770 -682
rect 696 -693 770 -687
rect 696 -707 703 -693
rect 762 -709 770 -693
rect 902 -697 910 -689
rect 867 -703 910 -697
rect 718 -748 727 -717
rect 867 -717 875 -703
rect 781 -748 789 -717
rect 718 -750 789 -748
rect 1348 -729 1356 -725
rect 1348 -730 1466 -729
rect 718 -751 790 -750
rect 718 -756 815 -751
rect 78 -773 338 -759
rect 781 -760 815 -756
rect 717 -784 766 -776
rect 233 -804 613 -790
rect 44 -839 518 -825
rect 343 -840 529 -839
rect 600 -835 613 -804
rect 695 -821 703 -799
rect 717 -793 727 -784
rect 758 -791 766 -784
rect 781 -792 789 -760
rect 804 -765 815 -760
rect 890 -763 900 -730
rect 1282 -734 1466 -730
rect 1282 -736 1356 -734
rect 1282 -750 1289 -736
rect 1348 -752 1356 -736
rect 1419 -735 1466 -734
rect 1419 -749 1426 -735
rect 804 -775 845 -765
rect 890 -772 1187 -763
rect 890 -798 900 -772
rect 1101 -773 1187 -772
rect 1179 -796 1187 -773
rect 1304 -791 1313 -760
rect 1367 -791 1375 -760
rect 1304 -793 1375 -791
rect 1482 -754 1489 -738
rect 1441 -790 1450 -759
rect 1499 -788 1507 -763
rect 1441 -793 1491 -790
rect 1304 -794 1376 -793
rect 1386 -794 1491 -793
rect 1179 -797 1267 -796
rect 1304 -797 1491 -794
rect 1499 -792 5056 -788
rect 1179 -804 1293 -797
rect 1304 -798 1466 -797
rect 1304 -799 1450 -798
rect 1367 -800 1450 -799
rect 1367 -802 1388 -800
rect 1179 -805 1267 -804
rect 1179 -807 1187 -805
rect 866 -825 875 -809
rect 866 -831 901 -825
rect 1303 -827 1352 -819
rect -281 -860 215 -858
rect -281 -862 352 -860
rect -282 -873 352 -862
rect 1281 -864 1289 -842
rect 1303 -836 1313 -827
rect 1344 -834 1352 -827
rect 1367 -825 1428 -816
rect 1454 -818 1462 -798
rect 1499 -805 1507 -792
rect 1367 -835 1375 -825
rect 1420 -834 1428 -825
rect 1440 -826 1466 -818
rect 1482 -824 1489 -814
rect 1440 -835 1450 -826
rect -281 -874 352 -873
rect -281 -876 215 -874
rect -281 -879 -252 -876
rect 337 -1029 352 -874
rect 762 -882 770 -877
rect 696 -888 770 -882
rect 696 -902 703 -888
rect 762 -904 770 -888
rect 902 -892 910 -884
rect 867 -898 910 -892
rect 718 -943 727 -912
rect 867 -912 875 -898
rect 781 -943 789 -912
rect 718 -945 789 -943
rect 1348 -919 1356 -915
rect 1348 -920 1466 -919
rect 718 -946 790 -945
rect 718 -951 815 -946
rect 781 -955 815 -951
rect 717 -979 766 -971
rect 695 -1016 703 -994
rect 717 -988 727 -979
rect 758 -986 766 -979
rect 781 -987 789 -955
rect 804 -960 815 -955
rect 890 -958 900 -925
rect 1282 -924 1466 -920
rect 1282 -926 1356 -924
rect 1282 -940 1289 -926
rect 1348 -942 1356 -926
rect 1419 -925 1466 -924
rect 1419 -939 1426 -925
rect 890 -959 927 -958
rect 1101 -959 1187 -953
rect 804 -970 845 -960
rect 890 -963 1187 -959
rect 890 -967 1142 -963
rect 890 -993 900 -967
rect 920 -968 1142 -967
rect 1179 -986 1187 -963
rect 1304 -981 1313 -950
rect 1367 -981 1375 -950
rect 1304 -983 1375 -981
rect 1482 -944 1489 -928
rect 1441 -980 1450 -949
rect 1499 -974 1507 -953
rect 1499 -978 5257 -974
rect 1441 -983 1491 -980
rect 1304 -984 1376 -983
rect 1386 -984 1491 -983
rect 1179 -987 1267 -986
rect 1304 -987 1491 -984
rect 1179 -994 1293 -987
rect 1304 -988 1466 -987
rect 1304 -989 1450 -988
rect 1367 -990 1450 -989
rect 1367 -992 1388 -990
rect 1179 -995 1267 -994
rect 1179 -997 1187 -995
rect 866 -1020 875 -1004
rect 1303 -1017 1352 -1009
rect 866 -1026 901 -1020
rect 337 -1030 620 -1029
rect 337 -1039 601 -1030
rect 1281 -1054 1289 -1032
rect 1303 -1026 1313 -1017
rect 1344 -1024 1352 -1017
rect 1367 -1015 1428 -1006
rect 1453 -1008 1461 -988
rect 1499 -995 1507 -978
rect 1367 -1025 1375 -1015
rect 1420 -1024 1428 -1015
rect 1440 -1016 1466 -1008
rect 1482 -1014 1489 -1004
rect 1440 -1025 1450 -1016
<< m2contact >>
rect 42 2370 70 2394
rect -282 903 -252 921
rect 207 2219 217 2232
rect 111 1727 135 1744
rect 132 1307 147 1322
rect 207 2108 215 2115
rect 388 2422 401 2435
rect 371 2219 381 2232
rect 372 2108 382 2116
rect 340 1804 351 1817
rect 322 1489 328 1496
rect 358 962 368 976
rect 286 512 303 521
rect 341 351 351 368
rect 45 67 68 74
<< metal2 >>
rect 185 2435 199 2436
rect 185 2423 388 2435
rect 185 2405 199 2423
rect 0 2394 199 2405
rect 0 2391 42 2394
rect 70 2391 199 2394
rect 43 1542 69 2370
rect 217 2219 371 2232
rect 215 2108 372 2115
rect 341 1744 351 1804
rect 135 1727 351 1744
rect -344 950 -328 952
rect -344 935 -342 950
rect -344 921 -328 935
rect -344 903 -282 921
rect 45 74 68 1542
rect 328 1489 329 1496
rect 322 1358 329 1489
rect 144 1357 330 1358
rect 133 1349 330 1357
rect 133 1322 148 1349
rect 147 1307 148 1322
rect 133 521 148 1307
rect 322 1001 329 1349
rect 132 512 286 521
rect 133 500 148 512
rect 341 368 351 1727
rect 357 962 358 976
rect 368 962 395 976
rect 341 349 351 351
rect 45 65 68 67
<< m3contact >>
rect -342 935 -328 950
rect 395 962 404 976
<< metal3 >>
rect 395 976 404 977
rect 395 950 404 962
rect -328 941 404 950
rect -328 935 403 941
<< labels >>
rlabel metal1 422 1666 423 1670 1 gnd
rlabel metal1 455 1791 456 1795 5 vdd
rlabel metal1 625 1666 626 1670 1 gnd
rlabel metal1 658 1791 659 1795 5 vdd
rlabel metal1 812 1666 813 1670 1 gnd
rlabel metal1 845 1791 846 1795 5 vdd
rlabel metal1 993 1666 994 1670 1 gnd
rlabel metal1 1026 1791 1027 1795 5 vdd
rlabel metal1 442 1349 443 1353 1 gnd
rlabel metal1 475 1474 476 1478 5 vdd
rlabel metal1 645 1349 646 1353 1 gnd
rlabel metal1 678 1474 679 1478 5 vdd
rlabel metal1 832 1349 833 1353 1 gnd
rlabel metal1 865 1474 866 1478 5 vdd
rlabel metal1 1013 1349 1014 1353 1 gnd
rlabel metal1 1046 1474 1047 1478 5 vdd
rlabel metal1 440 1058 441 1062 1 gnd
rlabel metal1 473 1183 474 1187 5 vdd
rlabel metal1 643 1058 644 1062 1 gnd
rlabel metal1 676 1183 677 1187 5 vdd
rlabel metal1 830 1058 831 1062 1 gnd
rlabel metal1 863 1183 864 1187 5 vdd
rlabel metal1 1011 1058 1012 1062 1 gnd
rlabel metal1 1044 1183 1045 1187 5 vdd
rlabel metal1 1398 1506 1399 1510 5 vdd
rlabel metal1 1365 1381 1366 1385 1 gnd
rlabel metal1 1535 1507 1536 1511 5 vdd
rlabel metal1 1629 1486 1632 1489 1 vdd
rlabel metal1 1629 1409 1633 1411 1 gnd
rlabel polysilicon 375 1837 377 1838 1 a1
rlabel polysilicon 411 1520 413 1521 1 a2
rlabel polysilicon 395 1230 397 1231 1 a3
rlabel polysilicon 374 1810 376 1811 1 b1
rlabel polycontact 390 1491 392 1492 1 b2
rlabel polycontact 388 1201 390 1202 1 b3
rlabel metal1 1142 1767 1145 1770 1 vdd
rlabel metal1 1142 1690 1146 1692 1 gnd
rlabel metal1 1167 1373 1171 1375 1 gnd
rlabel metal1 1167 1450 1170 1453 1 vdd
rlabel metal1 1176 1082 1180 1084 1 gnd
rlabel metal1 1176 1159 1179 1162 1 vdd
rlabel metal1 1140 1982 1144 1984 1 gnd
rlabel metal1 1140 2059 1143 2062 1 vdd
rlabel polysilicon 360 2098 362 2099 1 b0
rlabel polysilicon 367 2124 369 2125 1 a0
rlabel metal1 1020 2080 1021 2084 5 vdd
rlabel metal1 987 1955 988 1959 1 gnd
rlabel metal1 839 2080 840 2084 5 vdd
rlabel metal1 806 1955 807 1959 1 gnd
rlabel metal1 652 2080 653 2084 5 vdd
rlabel metal1 619 1955 620 1959 1 gnd
rlabel metal1 449 2080 450 2084 5 vdd
rlabel metal1 416 1955 417 1959 1 gnd
rlabel metal1 886 2344 888 2346 1 gnd
rlabel metal1 876 2473 878 2475 5 vdd
rlabel metal1 569 2470 570 2474 5 vdd
rlabel metal1 536 2345 537 2349 1 gnd
rlabel metal1 816 2564 818 2566 1 gnd
rlabel metal1 806 2693 808 2695 5 vdd
rlabel metal1 527 2564 528 2568 1 gnd
rlabel metal1 560 2689 561 2693 5 vdd
rlabel metal1 786 2854 788 2856 5 vdd
rlabel metal1 796 2725 798 2727 1 gnd
rlabel metal1 455 2609 458 2612 1 vdd
rlabel metal1 455 2532 459 2534 1 gnd
rlabel metal1 454 2849 458 2851 1 gnd
rlabel metal1 454 2926 457 2929 1 vdd
rlabel metal1 547 2723 548 2727 1 gnd
rlabel metal1 580 2848 581 2852 5 vdd
rlabel metal1 456 2764 459 2767 1 vdd
rlabel metal1 456 2687 460 2689 1 gnd
rlabel metal1 455 2300 459 2302 1 gnd
rlabel metal1 455 2377 458 2380 1 vdd
rlabel metal1 1673 2834 1674 2836 1 gnd
rlabel metal1 1673 2924 1674 2926 5 vdd
rlabel metal1 1650 2875 1651 2876 1 out
rlabel metal1 1510 2830 1511 2831 1 gnd
rlabel metal1 1511 2926 1512 2927 5 vdd
rlabel metal1 1679 1443 1681 1444 1 equal
rlabel metal1 731 3009 733 3011 5 vdd
rlabel metal1 741 2880 743 2882 1 gnd
rlabel metal1 580 3017 581 3021 5 vdd
rlabel metal1 547 2892 548 2896 1 gnd
rlabel metal1 1750 2879 1752 2880 1 agb
rlabel metal1 832 78 834 80 1 gnd
rlabel metal1 822 207 824 209 5 vdd
rlabel metal1 515 204 516 208 5 vdd
rlabel metal1 482 79 483 83 1 gnd
rlabel metal1 762 298 764 300 1 gnd
rlabel metal1 752 427 754 429 5 vdd
rlabel metal1 473 298 474 302 1 gnd
rlabel metal1 506 423 507 427 5 vdd
rlabel metal1 732 588 734 590 5 vdd
rlabel metal1 742 459 744 461 1 gnd
rlabel metal1 401 343 404 346 1 vdd
rlabel metal1 401 266 405 268 1 gnd
rlabel metal1 400 583 404 585 1 gnd
rlabel metal1 400 660 403 663 1 vdd
rlabel metal1 493 457 494 461 1 gnd
rlabel metal1 526 582 527 586 5 vdd
rlabel metal1 402 498 405 501 1 vdd
rlabel metal1 402 421 406 423 1 gnd
rlabel metal1 401 34 405 36 1 gnd
rlabel metal1 401 111 404 114 1 vdd
rlabel metal1 677 743 679 745 5 vdd
rlabel metal1 687 614 689 616 1 gnd
rlabel metal1 526 751 527 755 5 vdd
rlabel metal1 493 626 494 630 1 gnd
rlabel metal1 1571 660 1572 661 5 vdd
rlabel metal1 1570 564 1571 565 1 gnd
rlabel metal1 1733 658 1734 660 5 vdd
rlabel metal1 1733 568 1734 570 1 gnd
rlabel metal1 1038 3470 1039 3472 5 vdd
rlabel metal1 1038 3380 1039 3382 1 gnd
rlabel metal1 948 3376 949 3377 1 gnd
rlabel metal1 949 3472 950 3473 5 vdd
rlabel metal1 688 3357 689 3361 1 gnd
rlabel metal1 721 3482 722 3486 5 vdd
rlabel metal1 882 3345 884 3347 1 gnd
rlabel metal1 872 3474 874 3476 5 vdd
rlabel metal1 405 3361 406 3365 1 gnd
rlabel metal1 438 3486 439 3490 5 vdd
rlabel metal1 599 3349 601 3351 1 gnd
rlabel metal1 589 3478 591 3480 5 vdd
rlabel metal1 1849 3772 1850 3776 5 vdd
rlabel metal1 1816 3647 1817 3651 1 gnd
rlabel metal1 1668 3772 1669 3776 5 vdd
rlabel metal1 1635 3647 1636 3651 1 gnd
rlabel metal1 1481 3772 1482 3776 5 vdd
rlabel metal1 1448 3647 1449 3651 1 gnd
rlabel metal1 1278 3772 1279 3776 5 vdd
rlabel metal1 1245 3647 1246 3651 1 gnd
rlabel metal1 1109 3778 1110 3782 5 vdd
rlabel metal1 1076 3653 1077 3657 1 gnd
rlabel metal1 928 3778 929 3782 5 vdd
rlabel metal1 895 3653 896 3657 1 gnd
rlabel metal1 741 3778 742 3782 5 vdd
rlabel metal1 708 3653 709 3657 1 gnd
rlabel metal1 538 3778 539 3782 5 vdd
rlabel metal1 505 3653 506 3657 1 gnd
rlabel metal1 1010 4094 1011 4096 5 vdd
rlabel metal1 1010 4004 1011 4006 1 gnd
rlabel metal1 920 4000 921 4001 1 gnd
rlabel metal1 921 4096 922 4097 5 vdd
rlabel metal1 660 3981 661 3985 1 gnd
rlabel metal1 693 4106 694 4110 5 vdd
rlabel metal1 854 3969 856 3971 1 gnd
rlabel metal1 844 4098 846 4100 5 vdd
rlabel metal1 377 3985 378 3989 1 gnd
rlabel metal1 410 4110 411 4114 5 vdd
rlabel metal1 571 3973 573 3975 1 gnd
rlabel metal1 561 4102 563 4104 5 vdd
rlabel metal1 1821 4396 1822 4400 5 vdd
rlabel metal1 1788 4271 1789 4275 1 gnd
rlabel metal1 1640 4396 1641 4400 5 vdd
rlabel metal1 1607 4271 1608 4275 1 gnd
rlabel metal1 1453 4396 1454 4400 5 vdd
rlabel metal1 1420 4271 1421 4275 1 gnd
rlabel metal1 1250 4396 1251 4400 5 vdd
rlabel metal1 1217 4271 1218 4275 1 gnd
rlabel metal1 1081 4402 1082 4406 5 vdd
rlabel metal1 1048 4277 1049 4281 1 gnd
rlabel metal1 900 4402 901 4406 5 vdd
rlabel metal1 867 4277 868 4281 1 gnd
rlabel metal1 713 4402 714 4406 5 vdd
rlabel metal1 680 4277 681 4281 1 gnd
rlabel metal1 510 4402 511 4406 5 vdd
rlabel metal1 477 4277 478 4281 1 gnd
rlabel metal1 1030 4684 1031 4686 5 vdd
rlabel metal1 1030 4594 1031 4596 1 gnd
rlabel metal1 940 4590 941 4591 1 gnd
rlabel metal1 941 4686 942 4687 5 vdd
rlabel metal1 680 4571 681 4575 1 gnd
rlabel metal1 713 4696 714 4700 5 vdd
rlabel metal1 874 4559 876 4561 1 gnd
rlabel metal1 864 4688 866 4690 5 vdd
rlabel metal1 397 4575 398 4579 1 gnd
rlabel metal1 430 4700 431 4704 5 vdd
rlabel metal1 591 4563 593 4565 1 gnd
rlabel metal1 581 4692 583 4694 5 vdd
rlabel metal1 1841 4986 1842 4990 5 vdd
rlabel metal1 1808 4861 1809 4865 1 gnd
rlabel metal1 1660 4986 1661 4990 5 vdd
rlabel metal1 1627 4861 1628 4865 1 gnd
rlabel metal1 1473 4986 1474 4990 5 vdd
rlabel metal1 1440 4861 1441 4865 1 gnd
rlabel metal1 1270 4986 1271 4990 5 vdd
rlabel metal1 1237 4861 1238 4865 1 gnd
rlabel metal1 1101 4992 1102 4996 5 vdd
rlabel metal1 1068 4867 1069 4871 1 gnd
rlabel metal1 920 4992 921 4996 5 vdd
rlabel metal1 887 4867 888 4871 1 gnd
rlabel metal1 733 4992 734 4996 5 vdd
rlabel metal1 700 4867 701 4871 1 gnd
rlabel metal1 530 4992 531 4996 5 vdd
rlabel metal1 497 4867 498 4871 1 gnd
rlabel metal1 -626 4713 -625 4717 1 gnd
rlabel metal1 -593 4838 -592 4842 5 vdd
rlabel metal1 -423 4713 -422 4717 1 gnd
rlabel metal1 -390 4838 -389 4842 5 vdd
rlabel metal1 -236 4713 -235 4717 1 gnd
rlabel metal1 -203 4838 -202 4842 5 vdd
rlabel metal1 -55 4713 -54 4717 1 gnd
rlabel metal1 -22 4838 -21 4842 5 vdd
rlabel metal1 -626 5137 -625 5141 1 gnd
rlabel metal1 -593 5262 -592 5266 5 vdd
rlabel metal1 -423 5137 -422 5141 1 gnd
rlabel metal1 -390 5262 -389 5266 5 vdd
rlabel metal1 -236 5137 -235 5141 1 gnd
rlabel metal1 -203 5262 -202 5266 5 vdd
rlabel metal1 -55 5137 -54 5141 1 gnd
rlabel metal1 -22 5262 -21 5266 5 vdd
rlabel metal1 -626 5523 -625 5527 1 gnd
rlabel metal1 -593 5648 -592 5652 5 vdd
rlabel metal1 -423 5523 -422 5527 1 gnd
rlabel metal1 -390 5648 -389 5652 5 vdd
rlabel metal1 -236 5523 -235 5527 1 gnd
rlabel metal1 -203 5648 -202 5652 5 vdd
rlabel metal1 -55 5523 -54 5527 1 gnd
rlabel metal1 -22 5648 -21 5652 5 vdd
rlabel metal1 -50 5995 -49 5999 5 vdd
rlabel metal1 -83 5870 -82 5874 1 gnd
rlabel metal1 -231 5995 -230 5999 5 vdd
rlabel metal1 -264 5870 -263 5874 1 gnd
rlabel metal1 -418 5995 -417 5999 5 vdd
rlabel metal1 -451 5870 -450 5874 1 gnd
rlabel metal1 -621 5995 -620 5999 5 vdd
rlabel metal1 -654 5870 -653 5874 1 gnd
rlabel metal1 973 5408 974 5410 5 vdd
rlabel metal1 973 5318 974 5320 1 gnd
rlabel metal1 883 5314 884 5315 1 gnd
rlabel metal1 884 5410 885 5411 5 vdd
rlabel metal1 623 5295 624 5299 1 gnd
rlabel metal1 656 5420 657 5424 5 vdd
rlabel metal1 817 5283 819 5285 1 gnd
rlabel metal1 807 5412 809 5414 5 vdd
rlabel metal1 340 5299 341 5303 1 gnd
rlabel metal1 373 5424 374 5428 5 vdd
rlabel metal1 534 5287 536 5289 1 gnd
rlabel metal1 524 5416 526 5418 5 vdd
rlabel metal1 1784 5710 1785 5714 5 vdd
rlabel metal1 1751 5585 1752 5589 1 gnd
rlabel metal1 1603 5710 1604 5714 5 vdd
rlabel metal1 1570 5585 1571 5589 1 gnd
rlabel metal1 1416 5710 1417 5714 5 vdd
rlabel metal1 1383 5585 1384 5589 1 gnd
rlabel metal1 1213 5710 1214 5714 5 vdd
rlabel metal1 1180 5585 1181 5589 1 gnd
rlabel metal1 1044 5716 1045 5720 5 vdd
rlabel metal1 1011 5591 1012 5595 1 gnd
rlabel metal1 863 5716 864 5720 5 vdd
rlabel metal1 830 5591 831 5595 1 gnd
rlabel metal1 676 5716 677 5720 5 vdd
rlabel metal1 643 5591 644 5595 1 gnd
rlabel metal1 473 5716 474 5720 5 vdd
rlabel metal1 440 5591 441 5595 1 gnd
rlabel metal1 883 -304 885 -302 5 vdd
rlabel metal1 893 -433 895 -431 1 gnd
rlabel metal1 732 -296 733 -292 5 vdd
rlabel metal1 699 -421 700 -417 1 gnd
rlabel metal1 885 -502 887 -500 5 vdd
rlabel metal1 895 -631 897 -629 1 gnd
rlabel metal1 734 -494 735 -490 5 vdd
rlabel metal1 701 -619 702 -615 1 gnd
rlabel metal1 885 -700 887 -698 5 vdd
rlabel metal1 895 -829 897 -827 1 gnd
rlabel metal1 734 -692 735 -688 5 vdd
rlabel metal1 701 -817 702 -813 1 gnd
rlabel metal1 885 -895 887 -893 5 vdd
rlabel metal1 895 -1024 897 -1022 1 gnd
rlabel metal1 734 -887 735 -883 5 vdd
rlabel metal1 701 -1012 702 -1008 1 gnd
rlabel metal1 207 -439 210 -435 1 a0
rlabel metal1 231 -469 234 -465 1 b0
rlabel metal1 279 -494 282 -490 1 a1
rlabel metal1 261 -523 264 -519 1 b1
rlabel metal1 244 -764 247 -760 1 a2
rlabel metal1 279 -803 282 -799 1 b2
rlabel metal1 230 -834 233 -830 1 a3
rlabel metal1 215 -869 218 -865 1 b3
rlabel metal1 -1033 5943 -1027 5946 1 b0
rlabel metal1 -902 5672 -896 5675 1 b1
rlabel metal1 -930 5286 -924 5289 1 b2
rlabel metal1 -786 4865 -777 4867 1 b3
rlabel metal1 2380 5700 2382 5702 5 vdd
rlabel metal1 2390 5571 2392 5573 1 gnd
rlabel metal1 2229 5708 2230 5712 5 vdd
rlabel metal1 2196 5583 2197 5587 1 gnd
rlabel metal1 2378 4976 2380 4978 5 vdd
rlabel metal1 2388 4847 2390 4849 1 gnd
rlabel metal1 2227 4984 2228 4988 5 vdd
rlabel metal1 2194 4859 2195 4863 1 gnd
rlabel metal1 2379 4386 2381 4388 5 vdd
rlabel metal1 2389 4257 2391 4259 1 gnd
rlabel metal1 2228 4394 2229 4398 5 vdd
rlabel metal1 2195 4269 2196 4273 1 gnd
rlabel metal1 2196 3645 2197 3649 1 gnd
rlabel metal1 2229 3770 2230 3774 5 vdd
rlabel metal1 2390 3633 2392 3635 1 gnd
rlabel metal1 2380 3762 2382 3764 5 vdd
rlabel metal1 2198 3469 2199 3473 1 gnd
rlabel metal1 2231 3594 2232 3598 5 vdd
rlabel metal1 2392 3457 2394 3459 1 gnd
rlabel metal1 2382 3586 2384 3588 5 vdd
rlabel metal1 3034 5713 3037 5716 1 vdd
rlabel metal1 3034 5636 3038 5638 1 gnd
rlabel metal1 3161 5725 3163 5733 1 S1
rlabel metal1 3210 5721 3213 5725 1 S0
rlabel metal1 3305 5636 3308 5639 1 vdd
rlabel metal1 3305 5559 3309 5561 1 gnd
rlabel metal1 4671 852 4672 854 5 vdd
rlabel metal1 4671 762 4672 764 1 gnd
rlabel metal1 4549 758 4550 759 1 gnd
rlabel metal1 4550 854 4551 855 5 vdd
rlabel metal1 4915 1007 4916 1009 5 vdd
rlabel metal1 4915 917 4916 919 1 gnd
rlabel metal1 4793 913 4794 914 1 gnd
rlabel metal1 4794 1009 4795 1010 5 vdd
rlabel metal1 4688 807 4689 808 1 y0
rlabel metal1 4935 964 4936 965 1 y1
rlabel metal1 5172 1044 5173 1046 5 vdd
rlabel metal1 5172 954 5173 956 1 gnd
rlabel metal1 5050 950 5051 951 1 gnd
rlabel metal1 5051 1046 5052 1047 5 vdd
rlabel metal1 5192 1001 5193 1002 1 y2
rlabel metal1 5252 673 5253 674 5 vdd
rlabel metal1 5251 577 5252 578 1 gnd
rlabel metal1 5341 581 5342 583 1 gnd
rlabel metal1 5341 671 5342 673 5 vdd
rlabel metal1 5360 624 5362 626 1 y3
rlabel metal1 2405 3516 2407 3518 1 y4
rlabel metal1 2071 5648 2079 5650 1 ab0
rlabel metal1 2106 4925 2114 4927 1 ab1
rlabel metal1 2110 4334 2118 4336 1 ab2
rlabel metal1 2114 3709 2122 3711 1 ab3
rlabel metal1 2083 3671 2091 3673 1 ab4
rlabel metal1 1869 2740 1874 2746 1 co1
rlabel metal1 1928 1440 1933 1446 1 co2
rlabel space 1945 612 1950 618 1 co3
rlabel metal1 3360 5560 3361 5562 1 s0n
rlabel metal1 1483 -935 1486 -932 1 vdd
rlabel metal1 1483 -1012 1487 -1010 1 gnd
rlabel metal1 1457 -924 1458 -920 5 vdd
rlabel metal1 1287 -1050 1288 -1046 1 gnd
rlabel metal1 1320 -925 1321 -921 5 vdd
rlabel metal1 1320 -735 1321 -731 5 vdd
rlabel metal1 1287 -860 1288 -856 1 gnd
rlabel metal1 1457 -734 1458 -730 5 vdd
rlabel metal1 1483 -822 1487 -820 1 gnd
rlabel metal1 1483 -745 1486 -742 1 vdd
rlabel metal1 1483 -539 1486 -536 1 vdd
rlabel metal1 1483 -616 1487 -614 1 gnd
rlabel metal1 1457 -528 1458 -524 5 vdd
rlabel metal1 1287 -654 1288 -650 1 gnd
rlabel metal1 1320 -529 1321 -525 5 vdd
rlabel metal1 1320 -339 1321 -335 5 vdd
rlabel metal1 1287 -464 1288 -460 1 gnd
rlabel metal1 1457 -338 1458 -334 5 vdd
rlabel metal1 1483 -426 1487 -424 1 gnd
rlabel metal1 1483 -349 1486 -346 1 vdd
rlabel metal1 2282 668 2285 671 1 vdd
rlabel metal1 2282 591 2286 593 1 gnd
rlabel metal1 2256 679 2257 683 5 vdd
rlabel metal1 2086 553 2087 557 1 gnd
rlabel metal1 2119 678 2120 682 5 vdd
rlabel metal1 2119 1509 2120 1513 5 vdd
rlabel metal1 2086 1384 2087 1388 1 gnd
rlabel metal1 2256 1510 2257 1514 5 vdd
rlabel metal1 2282 1422 2286 1424 1 gnd
rlabel metal1 2282 1499 2285 1502 1 vdd
rlabel metal1 2119 2808 2120 2812 5 vdd
rlabel metal1 2086 2683 2087 2687 1 gnd
rlabel metal1 2256 2809 2257 2813 5 vdd
rlabel metal1 2282 2721 2286 2723 1 gnd
rlabel metal1 2282 2798 2285 2801 1 vdd
rlabel metal1 -1337 6251 -1331 6254 1 a1
rlabel metal1 -1423 6296 -1422 6298 1 a0
rlabel metal1 -1234 6193 -1228 6196 1 a2
rlabel metal1 -1222 6152 -1216 6155 1 a3
<< end >>
