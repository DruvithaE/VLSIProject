magic
tech scmos
timestamp 1700144367
<< nwell >>
rect 10 127 141 168
rect 213 127 344 168
rect 400 127 531 168
rect 581 127 712 168
rect 750 121 881 162
rect 953 121 1084 162
rect 1140 121 1271 162
rect 1321 121 1452 162
rect -90 -165 41 -124
rect 79 -176 145 -134
rect 193 -169 324 -128
rect 362 -180 428 -138
rect 457 -165 545 -140
rect 551 -165 604 -140
<< ntransistor >>
rect 36 57 43 72
rect 100 57 107 72
rect 239 57 246 72
rect 303 57 310 72
rect 426 57 435 72
rect 490 57 497 72
rect 607 57 614 72
rect 671 57 678 72
rect 776 51 783 66
rect 840 51 847 66
rect 979 51 986 66
rect 1043 51 1050 66
rect 1166 51 1173 66
rect 1230 51 1237 66
rect 1347 51 1354 66
rect 1411 51 1418 66
rect -64 -235 -57 -220
rect 0 -235 7 -220
rect 109 -241 117 -225
rect 219 -239 226 -224
rect 283 -239 290 -224
rect 479 -219 485 -208
rect 520 -219 526 -208
rect 571 -219 577 -208
rect 392 -245 400 -229
<< ptransistor >>
rect 36 142 43 157
rect 100 142 107 157
rect 239 142 246 157
rect 303 142 310 157
rect 426 142 433 157
rect 490 142 497 157
rect 607 142 614 157
rect 671 142 678 157
rect 776 136 783 151
rect 840 136 847 151
rect 979 136 986 151
rect 1043 136 1050 151
rect 1166 136 1173 151
rect 1230 136 1237 151
rect 1347 136 1354 151
rect 1411 136 1418 151
rect -64 -150 -57 -135
rect 0 -150 8 -135
rect 109 -163 117 -147
rect 219 -154 226 -139
rect 283 -154 290 -139
rect 392 -167 400 -151
rect 479 -158 485 -147
rect 520 -158 526 -147
rect 571 -158 577 -147
<< ndiffusion >>
rect 22 70 36 72
rect 22 63 24 70
rect 32 63 36 70
rect 22 57 36 63
rect 43 69 62 72
rect 43 60 46 69
rect 56 60 62 69
rect 43 57 62 60
rect 81 71 100 72
rect 81 63 87 71
rect 95 63 100 71
rect 81 57 100 63
rect 107 70 121 72
rect 107 62 110 70
rect 118 62 121 70
rect 107 57 121 62
rect 225 70 239 72
rect 225 63 227 70
rect 235 63 239 70
rect 225 57 239 63
rect 246 69 265 72
rect 246 60 249 69
rect 259 60 265 69
rect 246 57 265 60
rect 284 71 303 72
rect 284 63 290 71
rect 298 63 303 71
rect 284 57 303 63
rect 310 70 324 72
rect 310 62 313 70
rect 321 62 324 70
rect 310 57 324 62
rect 412 70 426 72
rect 412 63 414 70
rect 422 63 426 70
rect 412 57 426 63
rect 435 69 452 72
rect 435 60 436 69
rect 446 60 452 69
rect 435 57 452 60
rect 471 71 490 72
rect 471 63 477 71
rect 485 63 490 71
rect 471 57 490 63
rect 497 70 511 72
rect 497 62 500 70
rect 508 62 511 70
rect 497 57 511 62
rect 593 70 607 72
rect 593 63 595 70
rect 603 63 607 70
rect 593 57 607 63
rect 614 69 633 72
rect 614 60 617 69
rect 627 60 633 69
rect 614 57 633 60
rect 652 71 671 72
rect 652 63 658 71
rect 666 63 671 71
rect 652 57 671 63
rect 678 70 692 72
rect 678 62 681 70
rect 689 62 692 70
rect 678 57 692 62
rect 762 64 776 66
rect 762 57 764 64
rect 772 57 776 64
rect 762 51 776 57
rect 783 63 802 66
rect 783 54 786 63
rect 796 54 802 63
rect 783 51 802 54
rect 821 65 840 66
rect 821 57 827 65
rect 835 57 840 65
rect 821 51 840 57
rect 847 64 861 66
rect 847 56 850 64
rect 858 56 861 64
rect 847 51 861 56
rect 965 64 979 66
rect 965 57 967 64
rect 975 57 979 64
rect 965 51 979 57
rect 986 63 1005 66
rect 986 54 989 63
rect 999 54 1005 63
rect 986 51 1005 54
rect 1024 65 1043 66
rect 1024 57 1030 65
rect 1038 57 1043 65
rect 1024 51 1043 57
rect 1050 64 1064 66
rect 1050 56 1053 64
rect 1061 56 1064 64
rect 1050 51 1064 56
rect 1152 64 1166 66
rect 1152 57 1154 64
rect 1162 57 1166 64
rect 1152 51 1166 57
rect 1173 63 1192 66
rect 1173 54 1176 63
rect 1186 54 1192 63
rect 1173 51 1192 54
rect 1211 65 1230 66
rect 1211 57 1217 65
rect 1225 57 1230 65
rect 1211 51 1230 57
rect 1237 64 1251 66
rect 1237 56 1240 64
rect 1248 56 1251 64
rect 1237 51 1251 56
rect 1333 64 1347 66
rect 1333 57 1335 64
rect 1343 57 1347 64
rect 1333 51 1347 57
rect 1354 63 1373 66
rect 1354 54 1357 63
rect 1367 54 1373 63
rect 1354 51 1373 54
rect 1392 65 1411 66
rect 1392 57 1398 65
rect 1406 57 1411 65
rect 1392 51 1411 57
rect 1418 64 1432 66
rect 1418 56 1421 64
rect 1429 56 1432 64
rect 1418 51 1432 56
rect -78 -222 -64 -220
rect -78 -229 -76 -222
rect -68 -229 -64 -222
rect -78 -235 -64 -229
rect -57 -223 -38 -220
rect -57 -232 -54 -223
rect -44 -232 -38 -223
rect -57 -235 -38 -232
rect -19 -221 0 -220
rect -19 -229 -13 -221
rect -5 -229 0 -221
rect -19 -235 0 -229
rect 7 -222 21 -220
rect 7 -230 10 -222
rect 18 -230 21 -222
rect 7 -235 21 -230
rect 92 -229 109 -225
rect 92 -239 94 -229
rect 104 -239 109 -229
rect 92 -241 109 -239
rect 117 -228 132 -225
rect 117 -238 119 -228
rect 129 -238 132 -228
rect 117 -241 132 -238
rect 205 -226 219 -224
rect 205 -233 207 -226
rect 215 -233 219 -226
rect 205 -239 219 -233
rect 226 -227 245 -224
rect 226 -236 229 -227
rect 239 -236 245 -227
rect 226 -239 245 -236
rect 264 -225 283 -224
rect 264 -233 270 -225
rect 278 -233 283 -225
rect 264 -239 283 -233
rect 290 -226 304 -224
rect 290 -234 293 -226
rect 301 -234 304 -226
rect 468 -211 479 -208
rect 468 -216 470 -211
rect 476 -216 479 -211
rect 468 -219 479 -216
rect 485 -210 501 -208
rect 485 -216 489 -210
rect 496 -216 501 -210
rect 485 -219 501 -216
rect 506 -211 520 -208
rect 506 -216 510 -211
rect 516 -216 520 -211
rect 506 -219 520 -216
rect 526 -210 539 -208
rect 526 -216 529 -210
rect 536 -216 539 -210
rect 526 -219 539 -216
rect 555 -211 571 -208
rect 555 -216 561 -211
rect 567 -216 571 -211
rect 555 -219 571 -216
rect 577 -210 588 -208
rect 577 -216 579 -210
rect 586 -216 588 -210
rect 577 -219 588 -216
rect 290 -239 304 -234
rect 375 -233 392 -229
rect 375 -243 377 -233
rect 387 -243 392 -233
rect 375 -245 392 -243
rect 400 -232 415 -229
rect 400 -242 402 -232
rect 412 -242 415 -232
rect 400 -245 415 -242
<< pdiffusion >>
rect 22 155 36 157
rect 22 149 25 155
rect 32 149 36 155
rect 22 142 36 149
rect 43 153 62 157
rect 43 145 47 153
rect 56 145 62 153
rect 43 142 62 145
rect 89 153 100 157
rect 89 146 91 153
rect 99 146 100 153
rect 89 142 100 146
rect 107 151 129 157
rect 107 145 110 151
rect 118 145 129 151
rect 107 142 129 145
rect 225 155 239 157
rect 225 149 228 155
rect 235 149 239 155
rect 225 142 239 149
rect 246 153 265 157
rect 246 145 250 153
rect 259 145 265 153
rect 246 142 265 145
rect 292 153 303 157
rect 292 146 294 153
rect 302 146 303 153
rect 292 142 303 146
rect 310 151 332 157
rect 310 145 313 151
rect 321 145 332 151
rect 310 142 332 145
rect 412 155 426 157
rect 412 149 415 155
rect 422 149 426 155
rect 412 142 426 149
rect 433 153 452 157
rect 433 145 437 153
rect 446 145 452 153
rect 433 142 452 145
rect 479 153 490 157
rect 479 146 481 153
rect 489 146 490 153
rect 479 142 490 146
rect 497 151 519 157
rect 497 145 500 151
rect 508 145 519 151
rect 497 142 519 145
rect 593 155 607 157
rect 593 149 596 155
rect 603 149 607 155
rect 593 142 607 149
rect 614 153 633 157
rect 614 145 618 153
rect 627 145 633 153
rect 614 142 633 145
rect 660 153 671 157
rect 660 146 662 153
rect 670 146 671 153
rect 660 142 671 146
rect 678 151 700 157
rect 678 145 681 151
rect 689 145 700 151
rect 678 142 700 145
rect 762 149 776 151
rect 762 143 765 149
rect 772 143 776 149
rect 762 136 776 143
rect 783 147 802 151
rect 783 139 787 147
rect 796 139 802 147
rect 783 136 802 139
rect 829 147 840 151
rect 829 140 831 147
rect 839 140 840 147
rect 829 136 840 140
rect 847 145 869 151
rect 847 139 850 145
rect 858 139 869 145
rect 847 136 869 139
rect 965 149 979 151
rect 965 143 968 149
rect 975 143 979 149
rect 965 136 979 143
rect 986 147 1005 151
rect 986 139 990 147
rect 999 139 1005 147
rect 986 136 1005 139
rect 1032 147 1043 151
rect 1032 140 1034 147
rect 1042 140 1043 147
rect 1032 136 1043 140
rect 1050 145 1072 151
rect 1050 139 1053 145
rect 1061 139 1072 145
rect 1050 136 1072 139
rect 1152 149 1166 151
rect 1152 143 1155 149
rect 1162 143 1166 149
rect 1152 136 1166 143
rect 1173 147 1192 151
rect 1173 139 1177 147
rect 1186 139 1192 147
rect 1173 136 1192 139
rect 1219 147 1230 151
rect 1219 140 1221 147
rect 1229 140 1230 147
rect 1219 136 1230 140
rect 1237 145 1259 151
rect 1237 139 1240 145
rect 1248 139 1259 145
rect 1237 136 1259 139
rect 1333 149 1347 151
rect 1333 143 1336 149
rect 1343 143 1347 149
rect 1333 136 1347 143
rect 1354 147 1373 151
rect 1354 139 1358 147
rect 1367 139 1373 147
rect 1354 136 1373 139
rect 1400 147 1411 151
rect 1400 140 1402 147
rect 1410 140 1411 147
rect 1400 136 1411 140
rect 1418 145 1440 151
rect 1418 139 1421 145
rect 1429 139 1440 145
rect 1418 136 1440 139
rect -78 -137 -64 -135
rect -78 -143 -75 -137
rect -68 -143 -64 -137
rect -78 -150 -64 -143
rect -57 -139 -38 -135
rect -57 -147 -53 -139
rect -44 -147 -38 -139
rect -57 -150 -38 -147
rect -11 -139 0 -135
rect -11 -146 -9 -139
rect -1 -146 0 -139
rect -11 -150 0 -146
rect 8 -141 29 -135
rect 8 -147 10 -141
rect 18 -147 29 -141
rect 8 -150 29 -147
rect 93 -157 95 -147
rect 105 -157 109 -147
rect 93 -163 109 -157
rect 117 -150 133 -147
rect 117 -160 119 -150
rect 129 -160 133 -150
rect 117 -163 133 -160
rect 205 -141 219 -139
rect 205 -147 208 -141
rect 215 -147 219 -141
rect 205 -154 219 -147
rect 226 -143 245 -139
rect 226 -151 230 -143
rect 239 -151 245 -143
rect 226 -154 245 -151
rect 272 -143 283 -139
rect 272 -150 274 -143
rect 282 -150 283 -143
rect 272 -154 283 -150
rect 290 -145 312 -139
rect 290 -151 293 -145
rect 301 -151 312 -145
rect 468 -149 479 -147
rect 290 -154 312 -151
rect 376 -161 378 -151
rect 388 -161 392 -151
rect 376 -167 392 -161
rect 400 -154 416 -151
rect 400 -164 402 -154
rect 412 -164 416 -154
rect 468 -155 470 -149
rect 476 -155 479 -149
rect 468 -158 479 -155
rect 485 -152 501 -147
rect 485 -158 489 -152
rect 495 -158 501 -152
rect 506 -152 520 -147
rect 506 -158 510 -152
rect 516 -158 520 -152
rect 526 -152 539 -147
rect 526 -158 530 -152
rect 536 -158 539 -152
rect 558 -149 571 -147
rect 558 -155 561 -149
rect 567 -155 571 -149
rect 558 -158 571 -155
rect 577 -151 591 -147
rect 577 -157 579 -151
rect 586 -157 591 -151
rect 577 -158 591 -157
rect 400 -167 416 -164
<< ndcontact >>
rect 24 63 32 70
rect 46 60 56 69
rect 87 63 95 71
rect 110 62 118 70
rect 227 63 235 70
rect 249 60 259 69
rect 290 63 298 71
rect 313 62 321 70
rect 414 63 422 70
rect 436 60 446 69
rect 477 63 485 71
rect 500 62 508 70
rect 595 63 603 70
rect 617 60 627 69
rect 658 63 666 71
rect 681 62 689 70
rect 764 57 772 64
rect 786 54 796 63
rect 827 57 835 65
rect 850 56 858 64
rect 967 57 975 64
rect 989 54 999 63
rect 1030 57 1038 65
rect 1053 56 1061 64
rect 1154 57 1162 64
rect 1176 54 1186 63
rect 1217 57 1225 65
rect 1240 56 1248 64
rect 1335 57 1343 64
rect 1357 54 1367 63
rect 1398 57 1406 65
rect 1421 56 1429 64
rect -76 -229 -68 -222
rect -54 -232 -44 -223
rect -13 -229 -5 -221
rect 10 -230 18 -222
rect 94 -239 104 -229
rect 119 -238 129 -228
rect 207 -233 215 -226
rect 229 -236 239 -227
rect 270 -233 278 -225
rect 293 -234 301 -226
rect 470 -216 476 -211
rect 489 -216 496 -210
rect 510 -216 516 -211
rect 529 -216 536 -210
rect 561 -216 567 -211
rect 579 -216 586 -210
rect 377 -243 387 -233
rect 402 -242 412 -232
<< pdcontact >>
rect 25 149 32 155
rect 47 145 56 153
rect 91 146 99 153
rect 110 145 118 151
rect 228 149 235 155
rect 250 145 259 153
rect 294 146 302 153
rect 313 145 321 151
rect 415 149 422 155
rect 437 145 446 153
rect 481 146 489 153
rect 500 145 508 151
rect 596 149 603 155
rect 618 145 627 153
rect 662 146 670 153
rect 681 145 689 151
rect 765 143 772 149
rect 787 139 796 147
rect 831 140 839 147
rect 850 139 858 145
rect 968 143 975 149
rect 990 139 999 147
rect 1034 140 1042 147
rect 1053 139 1061 145
rect 1155 143 1162 149
rect 1177 139 1186 147
rect 1221 140 1229 147
rect 1240 139 1248 145
rect 1336 143 1343 149
rect 1358 139 1367 147
rect 1402 140 1410 147
rect 1421 139 1429 145
rect -75 -143 -68 -137
rect -53 -147 -44 -139
rect -9 -146 -1 -139
rect 10 -147 18 -141
rect 95 -157 105 -147
rect 119 -160 129 -150
rect 208 -147 215 -141
rect 230 -151 239 -143
rect 274 -150 282 -143
rect 293 -151 301 -145
rect 378 -161 388 -151
rect 402 -164 412 -154
rect 470 -155 476 -149
rect 489 -158 495 -152
rect 510 -158 516 -152
rect 530 -158 536 -152
rect 561 -155 567 -149
rect 579 -157 586 -151
<< polysilicon >>
rect 100 221 447 222
rect 108 214 447 221
rect 36 157 43 160
rect 100 157 107 210
rect 239 157 246 160
rect 303 157 310 160
rect 426 157 433 214
rect 840 208 855 216
rect 490 157 497 160
rect 607 157 614 190
rect 671 157 678 160
rect 776 151 783 154
rect 840 151 847 208
rect 1171 216 1627 218
rect 866 209 1627 216
rect 866 208 1187 209
rect 979 151 986 154
rect 1043 151 1050 154
rect 1166 151 1173 208
rect 1230 151 1237 154
rect 1347 151 1354 184
rect 1411 151 1418 154
rect 36 110 43 142
rect 36 72 43 99
rect 100 72 107 142
rect 239 72 246 142
rect 303 72 310 142
rect 426 76 433 142
rect 426 72 435 76
rect 490 72 497 142
rect 607 72 614 142
rect 671 72 678 142
rect 776 99 783 136
rect 776 66 783 90
rect 840 66 847 136
rect 979 66 986 136
rect 1043 66 1050 136
rect 1166 66 1173 136
rect 1230 66 1237 136
rect 1347 66 1354 136
rect 1411 66 1418 136
rect 36 13 43 57
rect 100 52 107 57
rect 239 13 246 57
rect 303 28 310 57
rect 36 6 246 13
rect 172 -50 186 6
rect 426 -34 435 57
rect 490 29 497 57
rect 607 53 614 57
rect 671 10 678 57
rect 776 7 783 51
rect 840 46 847 51
rect 979 7 986 51
rect 1043 22 1050 51
rect 1166 47 1173 51
rect 1230 23 1237 51
rect 1347 47 1354 51
rect 776 0 986 7
rect 1411 4 1418 51
rect 337 -44 443 -34
rect 1560 -41 1583 209
rect 173 -57 185 -50
rect -115 -74 47 -62
rect 183 -68 185 -57
rect 339 -60 346 -44
rect 426 -51 435 -44
rect 742 -57 1585 -41
rect 339 -74 346 -73
rect -115 -182 -103 -74
rect 743 -94 752 -57
rect 1560 -63 1583 -57
rect 0 -103 752 -94
rect -64 -135 -57 -132
rect 0 -135 8 -103
rect 283 -113 284 -107
rect 109 -147 117 -141
rect 219 -139 226 -136
rect 283 -139 290 -113
rect -64 -182 -57 -150
rect -115 -195 -57 -182
rect -64 -220 -57 -195
rect 0 -167 8 -150
rect 0 -220 7 -167
rect 109 -194 117 -163
rect 75 -195 117 -194
rect 85 -204 117 -195
rect 109 -225 117 -204
rect 174 -194 183 -142
rect 392 -151 400 -145
rect 479 -147 485 -143
rect 520 -147 526 -143
rect 571 -147 577 -143
rect 219 -193 226 -154
rect 190 -194 226 -193
rect 174 -202 226 -194
rect 136 -214 144 -204
rect 136 -219 145 -214
rect -64 -239 -57 -235
rect 0 -240 7 -235
rect 109 -249 117 -241
rect 136 -270 144 -219
rect 219 -224 226 -202
rect 283 -224 290 -154
rect 392 -198 400 -167
rect 358 -199 400 -198
rect 368 -208 400 -199
rect 479 -208 485 -158
rect 520 -208 526 -158
rect 571 -180 577 -158
rect 557 -186 577 -180
rect 571 -208 577 -186
rect 392 -229 400 -208
rect 219 -243 226 -239
rect 283 -244 290 -239
rect 392 -253 400 -245
rect 479 -269 485 -219
rect 432 -270 486 -269
rect 136 -276 486 -270
rect 137 -277 486 -276
rect 520 -294 526 -219
rect 571 -224 577 -219
rect 427 -295 526 -294
rect 439 -303 526 -295
rect 439 -304 521 -303
<< polycontact >>
rect 99 210 108 221
rect 607 190 614 197
rect 855 207 866 217
rect 1347 184 1354 191
rect 36 99 43 110
rect 775 90 784 99
rect 303 20 310 28
rect 490 21 497 29
rect 671 3 678 10
rect 1043 14 1050 22
rect 1230 15 1237 23
rect 1411 -3 1418 4
rect 47 -74 57 -59
rect 173 -68 183 -57
rect 339 -73 346 -60
rect 284 -113 290 -107
rect 173 -142 183 -131
rect 74 -205 85 -195
rect 136 -204 144 -192
rect 357 -209 368 -199
rect 552 -186 557 -180
rect 427 -307 439 -295
<< metal1 >>
rect -76 228 870 242
rect -76 210 99 221
rect -76 208 108 210
rect 854 217 867 228
rect 854 207 855 217
rect 866 207 867 217
rect 356 197 615 199
rect 79 186 341 196
rect 356 190 607 197
rect 614 190 615 197
rect 1096 191 1355 193
rect 356 189 615 190
rect -76 164 -12 176
rect 91 175 99 186
rect 294 175 302 186
rect -59 163 -12 164
rect -24 141 -12 163
rect 25 169 99 175
rect 25 155 32 169
rect 91 153 99 169
rect -21 113 -12 141
rect 228 169 302 175
rect 228 155 235 169
rect 47 114 56 145
rect 294 153 302 169
rect 110 124 118 145
rect 109 114 118 124
rect -21 110 43 113
rect -21 101 36 110
rect 47 111 118 114
rect 250 114 259 145
rect 313 114 321 145
rect 250 113 321 114
rect 357 113 366 189
rect 481 175 489 184
rect 662 175 670 184
rect 740 180 1081 190
rect 1096 184 1347 191
rect 1354 184 1355 191
rect 1096 183 1355 184
rect 415 169 489 175
rect 415 155 422 169
rect 481 153 489 169
rect 47 106 144 111
rect 250 106 366 113
rect 596 169 670 175
rect 831 169 839 180
rect 1034 169 1042 180
rect 596 155 603 169
rect 437 114 446 145
rect 662 153 670 169
rect 500 114 508 145
rect 437 113 508 114
rect 765 163 839 169
rect 618 114 627 145
rect 681 114 689 145
rect 765 149 772 163
rect 831 147 839 163
rect 618 113 689 114
rect 968 163 1042 169
rect 968 149 975 163
rect 437 106 554 113
rect 618 106 712 113
rect 110 102 144 106
rect 46 78 95 86
rect 24 41 32 63
rect 46 69 56 78
rect 87 71 95 78
rect 110 70 118 102
rect 133 29 144 102
rect 313 104 366 106
rect 500 104 554 106
rect 249 78 298 86
rect 227 41 235 63
rect 249 69 259 78
rect 290 71 298 78
rect 313 70 321 104
rect 436 78 485 86
rect 414 41 422 63
rect 436 69 446 78
rect 477 71 485 78
rect 500 70 508 104
rect 133 28 490 29
rect 133 20 303 28
rect 310 21 490 28
rect 497 21 531 29
rect 310 20 531 21
rect 133 18 531 20
rect 542 10 554 104
rect 681 104 712 106
rect 617 78 666 86
rect 595 41 603 63
rect 617 69 627 78
rect 658 71 666 78
rect 681 70 689 104
rect 704 98 712 104
rect 787 108 796 139
rect 1034 147 1042 163
rect 850 118 858 139
rect 849 108 858 118
rect 787 105 858 108
rect 990 108 999 139
rect 1053 108 1061 139
rect 990 107 1061 108
rect 1097 107 1106 183
rect 1221 169 1229 178
rect 1402 169 1410 178
rect 1155 163 1229 169
rect 1155 149 1162 163
rect 1221 147 1229 163
rect 787 100 884 105
rect 990 100 1106 107
rect 1336 163 1410 169
rect 1336 149 1343 163
rect 1177 108 1186 139
rect 1402 147 1410 163
rect 1240 108 1248 139
rect 1177 107 1248 108
rect 1358 108 1367 139
rect 1421 108 1429 139
rect 1358 107 1429 108
rect 1177 100 1294 107
rect 1358 100 1627 107
rect 704 90 775 98
rect 704 89 784 90
rect 850 96 884 100
rect 542 3 671 10
rect 678 3 711 10
rect 542 0 711 3
rect 726 -18 739 89
rect 786 72 835 80
rect 764 35 772 57
rect 786 63 796 72
rect 827 65 835 72
rect 850 64 858 96
rect 873 23 884 96
rect 1053 98 1106 100
rect 1240 98 1294 100
rect 989 72 1038 80
rect 967 35 975 57
rect 989 63 999 72
rect 1030 65 1038 72
rect 1053 64 1061 98
rect 1176 72 1225 80
rect 1154 35 1162 57
rect 1176 63 1186 72
rect 1217 65 1225 72
rect 1240 64 1248 98
rect 873 22 1230 23
rect 873 14 1043 22
rect 1050 15 1230 22
rect 1237 15 1271 23
rect 1050 14 1271 15
rect 873 12 1271 14
rect 1282 4 1294 98
rect 1421 99 1627 100
rect 1421 98 1440 99
rect 1357 72 1406 80
rect 1335 35 1343 57
rect 1357 63 1367 72
rect 1398 65 1406 72
rect 1421 64 1429 98
rect 1469 64 1627 67
rect 1468 53 1627 64
rect 1468 51 1491 53
rect 1547 51 1627 53
rect 1282 -3 1411 4
rect 1418 -3 1451 4
rect 1282 -6 1451 -3
rect 45 -30 742 -18
rect 48 -43 58 -30
rect 1468 -35 1484 51
rect 46 -59 58 -43
rect 1383 -48 1524 -35
rect 46 -73 47 -59
rect 57 -73 58 -59
rect -9 -117 -1 -112
rect -75 -123 -1 -117
rect -75 -137 -68 -123
rect -9 -139 -1 -123
rect 131 -127 139 -119
rect 96 -133 139 -127
rect 174 -131 183 -68
rect 339 -107 346 -73
rect 283 -113 284 -107
rect 290 -113 346 -107
rect 274 -121 282 -116
rect -53 -178 -44 -147
rect 96 -147 104 -133
rect 208 -127 282 -121
rect 208 -141 215 -127
rect 274 -143 282 -127
rect 414 -131 422 -123
rect 10 -178 18 -147
rect -53 -180 18 -178
rect -53 -181 19 -180
rect -53 -186 44 -181
rect 10 -190 44 -186
rect -54 -214 -5 -206
rect -76 -251 -68 -229
rect -54 -223 -44 -214
rect -13 -221 -5 -214
rect 10 -222 18 -190
rect 33 -195 44 -190
rect 119 -193 129 -160
rect 379 -137 422 -131
rect 230 -182 239 -151
rect 379 -151 387 -137
rect 470 -139 493 -133
rect 470 -149 476 -139
rect 293 -182 301 -151
rect 230 -184 301 -182
rect 561 -149 567 -133
rect 230 -185 302 -184
rect 230 -190 327 -185
rect 33 -205 74 -195
rect 119 -202 136 -193
rect 119 -228 129 -202
rect 144 -202 146 -193
rect 293 -194 327 -190
rect 229 -218 278 -210
rect 95 -255 104 -239
rect 207 -255 215 -233
rect 229 -227 239 -218
rect 270 -225 278 -218
rect 293 -226 301 -194
rect 316 -199 327 -194
rect 402 -197 412 -164
rect 489 -171 495 -158
rect 510 -171 516 -158
rect 489 -177 516 -171
rect 530 -180 536 -158
rect 579 -178 586 -157
rect 1383 -178 1392 -48
rect 530 -186 552 -180
rect 579 -186 1392 -178
rect 530 -192 536 -186
rect 316 -209 357 -199
rect 402 -205 440 -197
rect 489 -198 536 -192
rect 402 -206 439 -205
rect 402 -232 412 -206
rect 428 -212 439 -206
rect 489 -210 496 -198
rect 428 -217 440 -212
rect 529 -210 536 -198
rect 579 -187 1383 -186
rect 579 -210 586 -187
rect 95 -261 130 -255
rect 378 -259 387 -243
rect 378 -265 413 -259
rect 428 -295 439 -217
rect 470 -230 476 -216
rect 510 -230 516 -216
rect 470 -235 539 -230
rect 561 -233 567 -216
<< labels >>
rlabel metal1 30 45 31 49 1 gnd
rlabel metal1 63 170 64 174 5 vdd
rlabel metal1 233 45 234 49 1 gnd
rlabel metal1 266 170 267 174 5 vdd
rlabel metal1 420 45 421 49 1 gnd
rlabel metal1 453 170 454 174 5 vdd
rlabel metal1 601 45 602 49 1 gnd
rlabel metal1 634 170 635 174 5 vdd
rlabel metal1 770 39 771 43 1 gnd
rlabel metal1 803 164 804 168 5 vdd
rlabel metal1 973 39 974 43 1 gnd
rlabel metal1 1006 164 1007 168 5 vdd
rlabel metal1 1160 39 1161 43 1 gnd
rlabel metal1 1193 164 1194 168 5 vdd
rlabel metal1 1341 39 1342 43 1 gnd
rlabel metal1 1374 164 1375 168 5 vdd
rlabel metal1 114 -130 116 -128 5 vdd
rlabel metal1 124 -259 126 -257 1 gnd
rlabel metal1 -37 -122 -36 -118 5 vdd
rlabel metal1 -70 -247 -69 -243 1 gnd
rlabel metal1 397 -134 399 -132 5 vdd
rlabel metal1 407 -263 409 -261 1 gnd
rlabel metal1 246 -126 247 -122 5 vdd
rlabel metal1 213 -251 214 -247 1 gnd
rlabel metal1 474 -136 475 -135 5 vdd
rlabel metal1 473 -232 474 -231 1 gnd
rlabel metal1 563 -228 564 -226 1 gnd
rlabel metal1 563 -138 564 -136 5 vdd
<< end >>
