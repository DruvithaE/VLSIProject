magic
tech scmos
timestamp 1698574354
<< nwell >>
rect -187 -4 -121 38
rect -64 0 67 41
rect 139 0 270 41
rect 345 -1 549 41
<< ntransistor >>
rect -157 -69 -149 -53
rect -38 -70 -31 -55
rect 26 -70 33 -55
rect 165 -70 172 -55
rect 229 -70 236 -55
rect 376 -67 385 -52
rect 438 -67 447 -52
rect 500 -66 509 -51
<< ptransistor >>
rect -157 9 -149 25
rect -38 15 -31 30
rect 26 15 33 30
rect 165 15 172 30
rect 229 15 236 30
rect 376 13 385 28
rect 438 14 447 29
rect 500 13 509 28
<< ndiffusion >>
rect -174 -57 -157 -53
rect -174 -67 -172 -57
rect -162 -67 -157 -57
rect -174 -69 -157 -67
rect -149 -56 -134 -53
rect -149 -66 -147 -56
rect -137 -66 -134 -56
rect -149 -69 -134 -66
rect -52 -57 -38 -55
rect -52 -64 -50 -57
rect -42 -64 -38 -57
rect -52 -70 -38 -64
rect -31 -58 -12 -55
rect -31 -67 -28 -58
rect -18 -67 -12 -58
rect -31 -70 -12 -67
rect 7 -56 26 -55
rect 7 -64 13 -56
rect 21 -64 26 -56
rect 7 -70 26 -64
rect 33 -57 47 -55
rect 33 -65 36 -57
rect 44 -65 47 -57
rect 33 -70 47 -65
rect 151 -57 165 -55
rect 151 -64 153 -57
rect 161 -64 165 -57
rect 151 -70 165 -64
rect 172 -58 191 -55
rect 172 -67 175 -58
rect 185 -67 191 -58
rect 172 -70 191 -67
rect 210 -56 229 -55
rect 210 -64 216 -56
rect 224 -64 229 -56
rect 210 -70 229 -64
rect 236 -57 250 -55
rect 236 -65 239 -57
rect 247 -65 250 -57
rect 236 -70 250 -65
rect 363 -56 376 -52
rect 363 -65 364 -56
rect 374 -65 376 -56
rect 363 -67 376 -65
rect 385 -55 403 -52
rect 385 -64 387 -55
rect 397 -64 403 -55
rect 385 -67 403 -64
rect 423 -57 438 -52
rect 423 -66 425 -57
rect 435 -66 438 -57
rect 423 -67 438 -66
rect 447 -54 463 -52
rect 447 -63 450 -54
rect 460 -63 463 -54
rect 447 -67 463 -63
rect 485 -55 500 -51
rect 485 -64 488 -55
rect 498 -64 500 -55
rect 485 -66 500 -64
rect 509 -53 525 -51
rect 509 -62 513 -53
rect 523 -62 525 -53
rect 509 -66 525 -62
<< pdiffusion >>
rect -52 28 -38 30
rect -173 15 -171 25
rect -161 15 -157 25
rect -173 9 -157 15
rect -149 22 -133 25
rect -149 12 -147 22
rect -137 12 -133 22
rect -52 22 -49 28
rect -42 22 -38 28
rect -52 15 -38 22
rect -31 26 -12 30
rect -31 18 -27 26
rect -18 18 -12 26
rect -31 15 -12 18
rect 15 26 26 30
rect 15 19 17 26
rect 25 19 26 26
rect 15 15 26 19
rect 33 24 55 30
rect 33 18 36 24
rect 44 18 55 24
rect 33 15 55 18
rect 151 28 165 30
rect 151 22 154 28
rect 161 22 165 28
rect 151 15 165 22
rect 172 26 191 30
rect 172 18 176 26
rect 185 18 191 26
rect 172 15 191 18
rect 218 26 229 30
rect 218 19 220 26
rect 228 19 229 26
rect 218 15 229 19
rect 236 24 258 30
rect 236 18 239 24
rect 247 18 258 24
rect 236 15 258 18
rect 362 18 363 28
rect 374 18 376 28
rect -149 9 -133 12
rect 362 13 376 18
rect 385 23 402 28
rect 385 13 388 23
rect 398 13 402 23
rect 422 24 438 29
rect 422 16 426 24
rect 435 16 438 24
rect 422 14 438 16
rect 447 24 462 29
rect 447 15 450 24
rect 460 15 462 24
rect 447 14 462 15
rect 485 23 500 28
rect 485 14 488 23
rect 497 14 500 23
rect 485 13 500 14
rect 509 24 525 28
rect 509 15 513 24
rect 523 15 525 24
rect 509 13 525 15
<< ndcontact >>
rect -172 -67 -162 -57
rect -147 -66 -137 -56
rect -50 -64 -42 -57
rect -28 -67 -18 -58
rect 13 -64 21 -56
rect 36 -65 44 -57
rect 153 -64 161 -57
rect 175 -67 185 -58
rect 216 -64 224 -56
rect 239 -65 247 -57
rect 364 -65 374 -56
rect 387 -64 397 -55
rect 425 -66 435 -57
rect 450 -63 460 -54
rect 488 -64 498 -55
rect 513 -62 523 -53
<< pdcontact >>
rect -171 15 -161 25
rect -147 12 -137 22
rect -49 22 -42 28
rect -27 18 -18 26
rect 17 19 25 26
rect 36 18 44 24
rect 154 22 161 28
rect 176 18 185 26
rect 220 19 228 26
rect 239 18 247 24
rect 363 18 374 29
rect 388 13 398 23
rect 426 16 435 24
rect 450 15 460 24
rect 488 14 497 23
rect 513 15 523 24
<< polysilicon >>
rect -157 25 -149 31
rect -38 30 -31 33
rect 26 30 33 33
rect 165 30 172 33
rect 229 30 236 33
rect 376 28 385 35
rect 438 29 447 36
rect -157 -53 -149 9
rect -38 -55 -31 15
rect 26 -55 33 15
rect 165 -55 172 15
rect 229 -55 236 15
rect 500 28 509 36
rect 376 -13 385 13
rect 350 -23 385 -13
rect 376 -52 385 -23
rect 438 -52 447 14
rect 500 -51 509 13
rect -157 -77 -149 -69
rect -38 -74 -31 -70
rect 26 -75 33 -70
rect 165 -74 172 -70
rect 229 -75 236 -70
rect 376 -74 385 -67
rect 438 -98 447 -67
rect 500 -131 509 -66
<< polycontact >>
rect 338 -23 350 -13
rect 438 -111 448 -98
rect 500 -143 510 -131
<< metal1 >>
rect -135 59 403 69
rect -135 45 -127 59
rect 17 48 25 59
rect 220 48 228 59
rect -170 39 -127 45
rect -49 42 25 48
rect -170 25 -162 39
rect -49 28 -42 42
rect 17 26 25 42
rect -147 -21 -137 12
rect 154 42 228 48
rect 154 28 161 42
rect -27 -13 -18 18
rect 220 26 228 42
rect 364 43 375 59
rect 364 29 374 43
rect 36 -3 44 18
rect 35 -13 44 -3
rect -27 -16 44 -13
rect 176 -13 185 18
rect 239 -13 247 18
rect 388 -7 397 13
rect 426 -7 435 16
rect 176 -14 247 -13
rect -27 -21 70 -16
rect 176 -21 338 -14
rect -147 -30 -106 -21
rect -147 -56 -137 -30
rect -171 -83 -162 -67
rect -171 -89 -136 -83
rect -117 -131 -106 -30
rect 36 -25 70 -21
rect -28 -49 21 -41
rect -50 -86 -42 -64
rect -28 -58 -18 -49
rect 13 -56 21 -49
rect 36 -57 44 -25
rect 59 -98 70 -25
rect 239 -23 338 -21
rect 388 -17 435 -7
rect 451 -5 460 15
rect 488 -5 497 14
rect 451 -9 497 -5
rect 451 -15 496 -9
rect 513 -17 522 15
rect 175 -49 224 -41
rect 153 -86 161 -64
rect 175 -58 185 -49
rect 216 -56 224 -49
rect 239 -57 247 -23
rect 513 -26 538 -17
rect 513 -28 522 -26
rect 387 -38 522 -28
rect 388 -55 397 -38
rect 450 -54 459 -38
rect 513 -53 522 -38
rect 365 -79 374 -65
rect 426 -79 435 -66
rect 488 -79 497 -64
rect 364 -89 497 -79
rect 59 -109 438 -98
rect 344 -110 438 -109
rect -117 -143 500 -131
<< labels >>
rlabel polysilicon -35 -19 -34 -15 1 x
rlabel polysilicon 28 -29 29 -25 1 y
rlabel metal1 -44 -82 -43 -78 1 gnd
rlabel metal1 -11 43 -10 47 5 vdd
rlabel metal1 159 -82 160 -78 1 gnd
rlabel metal1 192 43 193 47 5 vdd
rlabel polysilicon -156 -27 -154 -25 1 z
rlabel metal1 -131 -26 -129 -24 1 zb
rlabel metal1 -152 42 -150 44 5 vdd
rlabel metal1 -142 -87 -140 -85 1 gnd
rlabel metal1 36 -20 39 -12 1 (x.y)b
rlabel polysilicon 166 -22 171 -7 1 a
rlabel polysilicon 230 -30 235 -15 1 b
rlabel metal1 242 -18 247 -13 1 (a.b)b
rlabel polysilicon 377 -23 380 -20 1 (a.b)b
rlabel polysilicon 441 -22 442 -18 1 (x.y)b
rlabel polysilicon 505 -22 506 -18 1 zb
rlabel metal1 366 49 368 53 1 vdd
rlabel metal1 370 -86 372 -81 1 gnd
rlabel metal1 525 -25 527 -20 1 finalout
<< end >>
