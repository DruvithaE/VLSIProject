magic
tech scmos
timestamp 1698587715
<< nwell >>
rect -53 0 167 25
<< ntransistor >>
rect -31 -54 -25 -43
rect 10 -54 16 -43
rect 49 -54 55 -43
rect 92 -54 98 -43
rect 134 -54 140 -43
<< ptransistor >>
rect -31 7 -25 18
rect 10 7 16 18
rect 49 7 55 18
rect 92 7 98 18
rect 134 7 140 18
<< ndiffusion >>
rect -42 -46 -31 -43
rect -42 -51 -40 -46
rect -34 -51 -31 -46
rect -42 -54 -31 -51
rect -25 -45 -9 -43
rect -25 -51 -21 -45
rect -14 -51 -9 -45
rect -25 -54 -9 -51
rect -4 -46 10 -43
rect -4 -51 0 -46
rect 6 -51 10 -46
rect -4 -54 10 -51
rect 16 -45 29 -43
rect 16 -51 19 -45
rect 26 -51 29 -45
rect 16 -54 29 -51
rect 35 -46 49 -43
rect 35 -52 39 -46
rect 45 -52 49 -46
rect 35 -54 49 -52
rect 55 -44 68 -43
rect 55 -51 58 -44
rect 65 -51 68 -44
rect 55 -54 68 -51
rect 78 -46 92 -43
rect 78 -52 82 -46
rect 88 -52 92 -46
rect 78 -54 92 -52
rect 98 -45 111 -43
rect 98 -51 100 -45
rect 107 -51 111 -45
rect 98 -54 111 -51
rect 118 -46 134 -43
rect 118 -51 124 -46
rect 130 -51 134 -46
rect 118 -54 134 -51
rect 140 -45 151 -43
rect 140 -51 142 -45
rect 149 -51 151 -45
rect 140 -54 151 -51
<< pdiffusion >>
rect -42 16 -31 18
rect -42 10 -40 16
rect -34 10 -31 16
rect -42 7 -31 10
rect -25 13 -9 18
rect -25 7 -21 13
rect -15 7 -9 13
rect -4 13 10 18
rect -4 7 0 13
rect 6 7 10 13
rect 16 13 29 18
rect 16 7 20 13
rect 26 7 29 13
rect 35 13 49 18
rect 35 7 39 13
rect 45 7 49 13
rect 55 13 68 18
rect 55 7 58 13
rect 64 7 68 13
rect 78 13 92 18
rect 78 7 82 13
rect 88 7 92 13
rect 98 13 111 18
rect 98 7 101 13
rect 107 7 111 13
rect 121 16 134 18
rect 121 10 124 16
rect 130 10 134 16
rect 121 7 134 10
rect 140 14 154 18
rect 140 8 142 14
rect 149 8 154 14
rect 140 7 154 8
<< ndcontact >>
rect -40 -51 -34 -46
rect -21 -51 -14 -45
rect 0 -51 6 -46
rect 19 -51 26 -45
rect 39 -52 45 -46
rect 58 -51 65 -44
rect 82 -52 88 -46
rect 100 -51 107 -45
rect 124 -51 130 -46
rect 142 -51 149 -45
<< pdcontact >>
rect -40 10 -34 16
rect -21 7 -15 13
rect 0 7 6 13
rect 20 7 26 13
rect 39 7 45 13
rect 58 7 64 13
rect 82 7 88 13
rect 101 7 107 13
rect 124 10 130 16
rect 142 8 149 14
<< polysilicon >>
rect -31 18 -25 22
rect 10 18 16 22
rect 49 18 55 22
rect 92 18 98 22
rect 134 18 140 22
rect -31 -43 -25 7
rect 10 -43 16 7
rect 49 -43 55 7
rect 92 -43 98 7
rect 134 -15 140 7
rect 120 -21 140 -15
rect 134 -43 140 -21
rect -31 -59 -25 -54
rect 10 -59 16 -54
rect 49 -59 55 -54
rect 92 -59 98 -54
rect 134 -59 140 -54
<< polycontact >>
rect 115 -21 120 -15
<< metal1 >>
rect -40 26 -17 32
rect -40 16 -34 26
rect 124 16 130 32
rect -21 -6 -15 7
rect 0 -6 6 7
rect -21 -12 6 -6
rect 20 -6 26 7
rect 39 -6 45 7
rect 20 -12 45 -6
rect 58 -6 64 7
rect 82 -6 88 7
rect 58 -12 88 -6
rect 101 -15 107 7
rect 142 -14 149 8
rect 101 -21 115 -15
rect 142 -20 156 -14
rect 101 -27 107 -21
rect -21 -33 107 -27
rect -21 -45 -14 -33
rect 19 -45 26 -33
rect 58 -44 65 -33
rect -40 -65 -34 -51
rect 0 -65 6 -51
rect 100 -45 107 -33
rect 39 -65 45 -52
rect 142 -45 149 -20
rect 82 -65 88 -52
rect -40 -70 88 -65
rect 124 -68 130 -51
<< labels >>
rlabel metal1 -36 29 -35 30 5 vdd
rlabel metal1 -37 -67 -36 -66 1 gnd
rlabel polysilicon -28 -18 -27 -17 1 a
rlabel polysilicon 13 -13 14 -12 1 b
rlabel polysilicon 51 -14 52 -13 1 c
rlabel polysilicon 94 -15 95 -14 1 d
rlabel metal1 103 -22 104 -21 1 out
rlabel metal1 126 27 127 29 5 vdd
rlabel metal1 126 -63 127 -61 1 gnd
rlabel metal1 142 -24 149 -7 1 fo
<< end >>
