magic
tech scmos
timestamp 1699701729
<< nwell >>
rect -14 0 33 25
<< ntransistor >>
rect 4 -43 10 -34
<< ptransistor >>
rect 4 8 10 17
<< ndiffusion >>
rect 2 -43 4 -34
rect 10 -43 12 -34
rect 20 -43 25 -34
<< pdiffusion >>
rect 2 8 4 17
rect 10 8 12 17
rect 21 8 25 17
<< ndcontact >>
rect -6 -43 2 -34
rect 12 -43 20 -34
<< pdcontact >>
rect -6 8 2 17
rect 12 8 21 17
<< polysilicon >>
rect 4 17 10 20
rect 4 -34 10 8
rect 4 -46 10 -43
<< metal1 >>
rect -5 17 2 33
rect 12 -34 20 8
rect -5 -53 2 -43
<< labels >>
rlabel metal1 -4 26 -1 29 1 vdd
rlabel metal1 -4 -51 0 -49 1 gnd
<< end >>
