magic
tech scmos
timestamp 1699877469
<< nwell >>
rect 10 127 141 168
rect 213 127 344 168
rect 400 127 531 168
rect 581 127 712 168
<< ntransistor >>
rect 36 57 43 72
rect 100 57 107 72
rect 239 57 246 72
rect 303 57 310 72
rect 426 57 433 72
rect 490 57 497 72
rect 607 57 614 72
rect 671 57 678 72
<< ptransistor >>
rect 36 142 43 157
rect 100 142 107 157
rect 239 142 246 157
rect 303 142 310 157
rect 426 142 433 157
rect 490 142 497 157
rect 607 142 614 157
rect 671 142 678 157
<< ndiffusion >>
rect 22 70 36 72
rect 22 63 24 70
rect 32 63 36 70
rect 22 57 36 63
rect 43 69 62 72
rect 43 60 46 69
rect 56 60 62 69
rect 43 57 62 60
rect 81 71 100 72
rect 81 63 87 71
rect 95 63 100 71
rect 81 57 100 63
rect 107 70 121 72
rect 107 62 110 70
rect 118 62 121 70
rect 107 57 121 62
rect 225 70 239 72
rect 225 63 227 70
rect 235 63 239 70
rect 225 57 239 63
rect 246 69 265 72
rect 246 60 249 69
rect 259 60 265 69
rect 246 57 265 60
rect 284 71 303 72
rect 284 63 290 71
rect 298 63 303 71
rect 284 57 303 63
rect 310 70 324 72
rect 310 62 313 70
rect 321 62 324 70
rect 310 57 324 62
rect 412 70 426 72
rect 412 63 414 70
rect 422 63 426 70
rect 412 57 426 63
rect 433 69 452 72
rect 433 60 436 69
rect 446 60 452 69
rect 433 57 452 60
rect 471 71 490 72
rect 471 63 477 71
rect 485 63 490 71
rect 471 57 490 63
rect 497 70 511 72
rect 497 62 500 70
rect 508 62 511 70
rect 497 57 511 62
rect 593 70 607 72
rect 593 63 595 70
rect 603 63 607 70
rect 593 57 607 63
rect 614 69 633 72
rect 614 60 617 69
rect 627 60 633 69
rect 614 57 633 60
rect 652 71 671 72
rect 652 63 658 71
rect 666 63 671 71
rect 652 57 671 63
rect 678 70 692 72
rect 678 62 681 70
rect 689 62 692 70
rect 678 57 692 62
<< pdiffusion >>
rect 22 155 36 157
rect 22 149 25 155
rect 32 149 36 155
rect 22 142 36 149
rect 43 153 62 157
rect 43 145 47 153
rect 56 145 62 153
rect 43 142 62 145
rect 89 153 100 157
rect 89 146 91 153
rect 99 146 100 153
rect 89 142 100 146
rect 107 151 129 157
rect 107 145 110 151
rect 118 145 129 151
rect 107 142 129 145
rect 225 155 239 157
rect 225 149 228 155
rect 235 149 239 155
rect 225 142 239 149
rect 246 153 265 157
rect 246 145 250 153
rect 259 145 265 153
rect 246 142 265 145
rect 292 153 303 157
rect 292 146 294 153
rect 302 146 303 153
rect 292 142 303 146
rect 310 151 332 157
rect 310 145 313 151
rect 321 145 332 151
rect 310 142 332 145
rect 412 155 426 157
rect 412 149 415 155
rect 422 149 426 155
rect 412 142 426 149
rect 433 153 452 157
rect 433 145 437 153
rect 446 145 452 153
rect 433 142 452 145
rect 479 153 490 157
rect 479 146 481 153
rect 489 146 490 153
rect 479 142 490 146
rect 497 151 519 157
rect 497 145 500 151
rect 508 145 519 151
rect 497 142 519 145
rect 593 155 607 157
rect 593 149 596 155
rect 603 149 607 155
rect 593 142 607 149
rect 614 153 633 157
rect 614 145 618 153
rect 627 145 633 153
rect 614 142 633 145
rect 660 153 671 157
rect 660 146 662 153
rect 670 146 671 153
rect 660 142 671 146
rect 678 151 700 157
rect 678 145 681 151
rect 689 145 700 151
rect 678 142 700 145
<< ndcontact >>
rect 24 63 32 70
rect 46 60 56 69
rect 87 63 95 71
rect 110 62 118 70
rect 227 63 235 70
rect 249 60 259 69
rect 290 63 298 71
rect 313 62 321 70
rect 414 63 422 70
rect 436 60 446 69
rect 477 63 485 71
rect 500 62 508 70
rect 595 63 603 70
rect 617 60 627 69
rect 658 63 666 71
rect 681 62 689 70
<< pdcontact >>
rect 25 149 32 155
rect 47 145 56 153
rect 91 146 99 153
rect 110 145 118 151
rect 228 149 235 155
rect 250 145 259 153
rect 294 146 302 153
rect 313 145 321 151
rect 415 149 422 155
rect 437 145 446 153
rect 481 146 489 153
rect 500 145 508 151
rect 596 149 603 155
rect 618 145 627 153
rect 662 146 670 153
rect 681 145 689 151
<< polysilicon >>
rect 100 214 447 222
rect 36 157 43 160
rect 100 157 107 214
rect 239 157 246 160
rect 303 157 310 160
rect 426 157 433 214
rect 490 157 497 160
rect 607 157 614 190
rect 671 157 678 160
rect 36 72 43 142
rect 100 72 107 142
rect 239 72 246 142
rect 303 72 310 142
rect 426 72 433 142
rect 490 72 497 142
rect 607 72 614 142
rect 671 72 678 142
rect 36 13 43 57
rect 100 52 107 57
rect 239 13 246 57
rect 303 28 310 57
rect 426 53 433 57
rect 490 29 497 57
rect 607 53 614 57
rect 36 6 246 13
rect 671 10 678 57
<< polycontact >>
rect 607 190 614 197
rect 303 20 310 28
rect 490 21 497 29
rect 671 3 678 10
<< metal1 >>
rect 356 197 615 199
rect 0 186 341 196
rect 356 190 607 197
rect 614 190 615 197
rect 356 189 615 190
rect 91 175 99 186
rect 294 175 302 186
rect 25 169 99 175
rect 25 155 32 169
rect 91 153 99 169
rect 228 169 302 175
rect 228 155 235 169
rect 47 114 56 145
rect 294 153 302 169
rect 110 124 118 145
rect 109 114 118 124
rect 47 111 118 114
rect 250 114 259 145
rect 313 114 321 145
rect 250 113 321 114
rect 357 113 366 189
rect 481 175 489 184
rect 662 175 670 184
rect 415 169 489 175
rect 415 155 422 169
rect 481 153 489 169
rect 47 106 144 111
rect 250 106 366 113
rect 596 169 670 175
rect 596 155 603 169
rect 437 114 446 145
rect 662 153 670 169
rect 500 114 508 145
rect 437 113 508 114
rect 618 114 627 145
rect 681 114 689 145
rect 618 113 689 114
rect 437 106 554 113
rect 618 106 709 113
rect 110 102 144 106
rect 46 78 95 86
rect 24 41 32 63
rect 46 69 56 78
rect 87 71 95 78
rect 110 70 118 102
rect 133 29 144 102
rect 313 104 366 106
rect 500 104 554 106
rect 249 78 298 86
rect 227 41 235 63
rect 249 69 259 78
rect 290 71 298 78
rect 313 70 321 104
rect 436 78 485 86
rect 414 41 422 63
rect 436 69 446 78
rect 477 71 485 78
rect 500 70 508 104
rect 133 28 490 29
rect 133 20 303 28
rect 310 21 490 28
rect 497 21 531 29
rect 310 20 531 21
rect 133 18 531 20
rect 542 10 554 104
rect 681 104 709 106
rect 617 78 666 86
rect 595 41 603 63
rect 617 69 627 78
rect 658 71 666 78
rect 681 70 689 104
rect 542 3 671 10
rect 678 3 711 10
rect 542 0 711 3
<< labels >>
rlabel metal1 30 45 31 49 1 gnd
rlabel metal1 63 170 64 174 5 vdd
rlabel metal1 233 45 234 49 1 gnd
rlabel metal1 266 170 267 174 5 vdd
rlabel metal1 420 45 421 49 1 gnd
rlabel metal1 453 170 454 174 5 vdd
rlabel metal1 601 45 602 49 1 gnd
rlabel metal1 634 170 635 174 5 vdd
<< end >>
