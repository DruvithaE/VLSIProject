magic
tech scmos
timestamp 1700166582
<< nwell >>
rect 41 1070 172 1111
rect 244 1070 375 1111
rect 431 1070 562 1111
rect 612 1070 743 1111
rect 47 735 178 776
rect 250 735 381 776
rect 437 735 568 776
rect 618 735 749 776
rect 67 418 198 459
rect 270 418 401 459
rect 457 418 588 459
rect 638 418 769 459
rect 990 450 1121 491
rect 1127 451 1258 492
rect 1978 186 2109 227
rect 2115 187 2246 228
rect 2282 189 2329 214
rect 65 127 196 168
rect 268 127 399 168
rect 455 127 586 168
rect 636 127 767 168
<< ntransistor >>
rect 67 1000 74 1015
rect 131 1000 138 1015
rect 270 1000 277 1015
rect 334 1000 341 1015
rect 457 1000 464 1015
rect 521 1000 528 1015
rect 638 1000 645 1015
rect 702 1000 709 1015
rect 73 665 80 680
rect 137 665 144 680
rect 276 665 283 680
rect 340 665 347 680
rect 463 665 470 680
rect 527 665 534 680
rect 644 665 651 680
rect 708 665 715 680
rect 1016 380 1023 395
rect 1080 380 1087 395
rect 1153 381 1160 396
rect 1217 381 1224 396
rect 93 348 100 363
rect 157 348 164 363
rect 296 348 303 363
rect 360 348 367 363
rect 483 348 490 363
rect 547 348 554 363
rect 664 348 671 363
rect 728 348 735 363
rect 2300 146 2306 155
rect 2004 116 2011 131
rect 2068 116 2075 131
rect 2141 117 2148 132
rect 2205 117 2212 132
rect 91 57 98 72
rect 155 57 162 72
rect 294 57 301 72
rect 358 57 365 72
rect 481 57 488 72
rect 545 57 552 72
rect 662 57 669 72
rect 726 57 733 72
<< ptransistor >>
rect 67 1085 74 1100
rect 131 1085 138 1100
rect 270 1085 277 1100
rect 334 1085 341 1100
rect 457 1085 464 1100
rect 521 1085 528 1100
rect 638 1085 645 1100
rect 702 1085 709 1100
rect 73 750 80 765
rect 137 750 144 765
rect 276 750 283 765
rect 340 750 347 765
rect 463 750 470 765
rect 527 750 534 765
rect 644 750 651 765
rect 708 750 715 765
rect 1016 465 1023 480
rect 1080 465 1087 480
rect 1153 466 1160 481
rect 1217 466 1224 481
rect 93 433 100 448
rect 157 433 164 448
rect 296 433 303 448
rect 360 433 367 448
rect 483 433 490 448
rect 547 433 554 448
rect 664 433 671 448
rect 728 433 735 448
rect 91 142 98 157
rect 155 142 162 157
rect 294 142 301 157
rect 358 142 365 157
rect 481 142 488 157
rect 545 142 552 157
rect 662 142 669 157
rect 726 142 733 157
rect 2004 201 2011 216
rect 2068 201 2075 216
rect 2141 202 2148 217
rect 2205 202 2212 217
rect 2300 197 2306 206
<< ndiffusion >>
rect 53 1013 67 1015
rect 53 1006 55 1013
rect 63 1006 67 1013
rect 53 1000 67 1006
rect 74 1012 93 1015
rect 74 1003 77 1012
rect 87 1003 93 1012
rect 74 1000 93 1003
rect 112 1014 131 1015
rect 112 1006 118 1014
rect 126 1006 131 1014
rect 112 1000 131 1006
rect 138 1013 152 1015
rect 138 1005 141 1013
rect 149 1005 152 1013
rect 138 1000 152 1005
rect 256 1013 270 1015
rect 256 1006 258 1013
rect 266 1006 270 1013
rect 256 1000 270 1006
rect 277 1012 296 1015
rect 277 1003 280 1012
rect 290 1003 296 1012
rect 277 1000 296 1003
rect 315 1014 334 1015
rect 315 1006 321 1014
rect 329 1006 334 1014
rect 315 1000 334 1006
rect 341 1013 355 1015
rect 341 1005 344 1013
rect 352 1005 355 1013
rect 341 1000 355 1005
rect 443 1013 457 1015
rect 443 1006 445 1013
rect 453 1006 457 1013
rect 443 1000 457 1006
rect 464 1012 483 1015
rect 464 1003 467 1012
rect 477 1003 483 1012
rect 464 1000 483 1003
rect 502 1014 521 1015
rect 502 1006 508 1014
rect 516 1006 521 1014
rect 502 1000 521 1006
rect 528 1013 542 1015
rect 528 1005 531 1013
rect 539 1005 542 1013
rect 528 1000 542 1005
rect 624 1013 638 1015
rect 624 1006 626 1013
rect 634 1006 638 1013
rect 624 1000 638 1006
rect 645 1012 664 1015
rect 645 1003 648 1012
rect 658 1003 664 1012
rect 645 1000 664 1003
rect 683 1014 702 1015
rect 683 1006 689 1014
rect 697 1006 702 1014
rect 683 1000 702 1006
rect 709 1013 723 1015
rect 709 1005 712 1013
rect 720 1005 723 1013
rect 709 1000 723 1005
rect 59 678 73 680
rect 59 671 61 678
rect 69 671 73 678
rect 59 665 73 671
rect 80 677 99 680
rect 80 668 83 677
rect 93 668 99 677
rect 80 665 99 668
rect 118 679 137 680
rect 118 671 124 679
rect 132 671 137 679
rect 118 665 137 671
rect 144 678 158 680
rect 144 670 147 678
rect 155 670 158 678
rect 144 665 158 670
rect 262 678 276 680
rect 262 671 264 678
rect 272 671 276 678
rect 262 665 276 671
rect 283 677 302 680
rect 283 668 286 677
rect 296 668 302 677
rect 283 665 302 668
rect 321 679 340 680
rect 321 671 327 679
rect 335 671 340 679
rect 321 665 340 671
rect 347 678 361 680
rect 347 670 350 678
rect 358 670 361 678
rect 347 665 361 670
rect 449 678 463 680
rect 449 671 451 678
rect 459 671 463 678
rect 449 665 463 671
rect 470 677 489 680
rect 470 668 473 677
rect 483 668 489 677
rect 470 665 489 668
rect 508 679 527 680
rect 508 671 514 679
rect 522 671 527 679
rect 508 665 527 671
rect 534 678 548 680
rect 534 670 537 678
rect 545 670 548 678
rect 534 665 548 670
rect 630 678 644 680
rect 630 671 632 678
rect 640 671 644 678
rect 630 665 644 671
rect 651 677 670 680
rect 651 668 654 677
rect 664 668 670 677
rect 651 665 670 668
rect 689 679 708 680
rect 689 671 695 679
rect 703 671 708 679
rect 689 665 708 671
rect 715 678 729 680
rect 715 670 718 678
rect 726 670 729 678
rect 715 665 729 670
rect 1002 393 1016 395
rect 1002 386 1004 393
rect 1012 386 1016 393
rect 1002 380 1016 386
rect 1023 392 1042 395
rect 1023 383 1026 392
rect 1036 383 1042 392
rect 1023 380 1042 383
rect 1061 394 1080 395
rect 1061 386 1067 394
rect 1075 386 1080 394
rect 1061 380 1080 386
rect 1087 393 1101 395
rect 1087 385 1090 393
rect 1098 385 1101 393
rect 1087 380 1101 385
rect 1137 394 1153 396
rect 1137 386 1143 394
rect 1151 386 1153 394
rect 1137 381 1153 386
rect 1160 393 1179 396
rect 1160 384 1163 393
rect 1173 384 1179 393
rect 1160 381 1179 384
rect 1198 395 1217 396
rect 1198 387 1204 395
rect 1212 387 1217 395
rect 1198 381 1217 387
rect 1224 394 1238 396
rect 1224 386 1227 394
rect 1235 386 1238 394
rect 1224 381 1238 386
rect 79 361 93 363
rect 79 354 81 361
rect 89 354 93 361
rect 79 348 93 354
rect 100 360 119 363
rect 100 351 103 360
rect 113 351 119 360
rect 100 348 119 351
rect 138 362 157 363
rect 138 354 144 362
rect 152 354 157 362
rect 138 348 157 354
rect 164 361 178 363
rect 164 353 167 361
rect 175 353 178 361
rect 164 348 178 353
rect 282 361 296 363
rect 282 354 284 361
rect 292 354 296 361
rect 282 348 296 354
rect 303 360 322 363
rect 303 351 306 360
rect 316 351 322 360
rect 303 348 322 351
rect 341 362 360 363
rect 341 354 347 362
rect 355 354 360 362
rect 341 348 360 354
rect 367 361 381 363
rect 367 353 370 361
rect 378 353 381 361
rect 367 348 381 353
rect 469 361 483 363
rect 469 354 471 361
rect 479 354 483 361
rect 469 348 483 354
rect 490 360 509 363
rect 490 351 493 360
rect 503 351 509 360
rect 490 348 509 351
rect 528 362 547 363
rect 528 354 534 362
rect 542 354 547 362
rect 528 348 547 354
rect 554 361 568 363
rect 554 353 557 361
rect 565 353 568 361
rect 554 348 568 353
rect 650 361 664 363
rect 650 354 652 361
rect 660 354 664 361
rect 650 348 664 354
rect 671 360 690 363
rect 671 351 674 360
rect 684 351 690 360
rect 671 348 690 351
rect 709 362 728 363
rect 709 354 715 362
rect 723 354 728 362
rect 709 348 728 354
rect 735 361 749 363
rect 735 353 738 361
rect 746 353 749 361
rect 735 348 749 353
rect 2298 146 2300 155
rect 2306 146 2308 155
rect 2316 146 2321 155
rect 1990 129 2004 131
rect 1990 122 1992 129
rect 2000 122 2004 129
rect 1990 116 2004 122
rect 2011 128 2030 131
rect 2011 119 2014 128
rect 2024 119 2030 128
rect 2011 116 2030 119
rect 2049 130 2068 131
rect 2049 122 2055 130
rect 2063 122 2068 130
rect 2049 116 2068 122
rect 2075 129 2089 131
rect 2075 121 2078 129
rect 2086 121 2089 129
rect 2075 116 2089 121
rect 2125 130 2141 132
rect 2125 122 2131 130
rect 2139 122 2141 130
rect 2125 117 2141 122
rect 2148 129 2167 132
rect 2148 120 2151 129
rect 2161 120 2167 129
rect 2148 117 2167 120
rect 2186 131 2205 132
rect 2186 123 2192 131
rect 2200 123 2205 131
rect 2186 117 2205 123
rect 2212 130 2226 132
rect 2212 122 2215 130
rect 2223 122 2226 130
rect 2212 117 2226 122
rect 77 70 91 72
rect 77 63 79 70
rect 87 63 91 70
rect 77 57 91 63
rect 98 69 117 72
rect 98 60 101 69
rect 111 60 117 69
rect 98 57 117 60
rect 136 71 155 72
rect 136 63 142 71
rect 150 63 155 71
rect 136 57 155 63
rect 162 70 176 72
rect 162 62 165 70
rect 173 62 176 70
rect 162 57 176 62
rect 280 70 294 72
rect 280 63 282 70
rect 290 63 294 70
rect 280 57 294 63
rect 301 69 320 72
rect 301 60 304 69
rect 314 60 320 69
rect 301 57 320 60
rect 339 71 358 72
rect 339 63 345 71
rect 353 63 358 71
rect 339 57 358 63
rect 365 70 379 72
rect 365 62 368 70
rect 376 62 379 70
rect 365 57 379 62
rect 467 70 481 72
rect 467 63 469 70
rect 477 63 481 70
rect 467 57 481 63
rect 488 69 507 72
rect 488 60 491 69
rect 501 60 507 69
rect 488 57 507 60
rect 526 71 545 72
rect 526 63 532 71
rect 540 63 545 71
rect 526 57 545 63
rect 552 70 566 72
rect 552 62 555 70
rect 563 62 566 70
rect 552 57 566 62
rect 648 70 662 72
rect 648 63 650 70
rect 658 63 662 70
rect 648 57 662 63
rect 669 69 688 72
rect 669 60 672 69
rect 682 60 688 69
rect 669 57 688 60
rect 707 71 726 72
rect 707 63 713 71
rect 721 63 726 71
rect 707 57 726 63
rect 733 70 747 72
rect 733 62 736 70
rect 744 62 747 70
rect 733 57 747 62
<< pdiffusion >>
rect 53 1098 67 1100
rect 53 1092 56 1098
rect 63 1092 67 1098
rect 53 1085 67 1092
rect 74 1096 93 1100
rect 74 1088 78 1096
rect 87 1088 93 1096
rect 74 1085 93 1088
rect 120 1096 131 1100
rect 120 1089 122 1096
rect 130 1089 131 1096
rect 120 1085 131 1089
rect 138 1094 160 1100
rect 138 1088 141 1094
rect 149 1088 160 1094
rect 138 1085 160 1088
rect 256 1098 270 1100
rect 256 1092 259 1098
rect 266 1092 270 1098
rect 256 1085 270 1092
rect 277 1096 296 1100
rect 277 1088 281 1096
rect 290 1088 296 1096
rect 277 1085 296 1088
rect 323 1096 334 1100
rect 323 1089 325 1096
rect 333 1089 334 1096
rect 323 1085 334 1089
rect 341 1094 363 1100
rect 341 1088 344 1094
rect 352 1088 363 1094
rect 341 1085 363 1088
rect 443 1098 457 1100
rect 443 1092 446 1098
rect 453 1092 457 1098
rect 443 1085 457 1092
rect 464 1096 483 1100
rect 464 1088 468 1096
rect 477 1088 483 1096
rect 464 1085 483 1088
rect 510 1096 521 1100
rect 510 1089 512 1096
rect 520 1089 521 1096
rect 510 1085 521 1089
rect 528 1094 550 1100
rect 528 1088 531 1094
rect 539 1088 550 1094
rect 528 1085 550 1088
rect 624 1098 638 1100
rect 624 1092 627 1098
rect 634 1092 638 1098
rect 624 1085 638 1092
rect 645 1096 664 1100
rect 645 1088 649 1096
rect 658 1088 664 1096
rect 645 1085 664 1088
rect 691 1096 702 1100
rect 691 1089 693 1096
rect 701 1089 702 1096
rect 691 1085 702 1089
rect 709 1094 731 1100
rect 709 1088 712 1094
rect 720 1088 731 1094
rect 709 1085 731 1088
rect 59 763 73 765
rect 59 757 62 763
rect 69 757 73 763
rect 59 750 73 757
rect 80 761 99 765
rect 80 753 84 761
rect 93 753 99 761
rect 80 750 99 753
rect 126 761 137 765
rect 126 754 128 761
rect 136 754 137 761
rect 126 750 137 754
rect 144 759 166 765
rect 144 753 147 759
rect 155 753 166 759
rect 144 750 166 753
rect 262 763 276 765
rect 262 757 265 763
rect 272 757 276 763
rect 262 750 276 757
rect 283 761 302 765
rect 283 753 287 761
rect 296 753 302 761
rect 283 750 302 753
rect 329 761 340 765
rect 329 754 331 761
rect 339 754 340 761
rect 329 750 340 754
rect 347 759 369 765
rect 347 753 350 759
rect 358 753 369 759
rect 347 750 369 753
rect 449 763 463 765
rect 449 757 452 763
rect 459 757 463 763
rect 449 750 463 757
rect 470 761 489 765
rect 470 753 474 761
rect 483 753 489 761
rect 470 750 489 753
rect 516 761 527 765
rect 516 754 518 761
rect 526 754 527 761
rect 516 750 527 754
rect 534 759 556 765
rect 534 753 537 759
rect 545 753 556 759
rect 534 750 556 753
rect 630 763 644 765
rect 630 757 633 763
rect 640 757 644 763
rect 630 750 644 757
rect 651 761 670 765
rect 651 753 655 761
rect 664 753 670 761
rect 651 750 670 753
rect 697 761 708 765
rect 697 754 699 761
rect 707 754 708 761
rect 697 750 708 754
rect 715 759 737 765
rect 715 753 718 759
rect 726 753 737 759
rect 715 750 737 753
rect 1002 478 1016 480
rect 1002 472 1005 478
rect 1012 472 1016 478
rect 1002 465 1016 472
rect 1023 476 1042 480
rect 1023 468 1027 476
rect 1036 468 1042 476
rect 1023 465 1042 468
rect 1069 476 1080 480
rect 1069 469 1071 476
rect 1079 469 1080 476
rect 1069 465 1080 469
rect 1087 474 1109 480
rect 1087 468 1090 474
rect 1098 468 1109 474
rect 1087 465 1109 468
rect 1139 479 1153 481
rect 1139 473 1142 479
rect 1149 473 1153 479
rect 1139 466 1153 473
rect 1160 477 1179 481
rect 1160 469 1164 477
rect 1173 469 1179 477
rect 1160 466 1179 469
rect 1206 477 1217 481
rect 1206 470 1208 477
rect 1216 470 1217 477
rect 1206 466 1217 470
rect 1224 475 1246 481
rect 1224 469 1227 475
rect 1235 469 1246 475
rect 1224 466 1246 469
rect 79 446 93 448
rect 79 440 82 446
rect 89 440 93 446
rect 79 433 93 440
rect 100 444 119 448
rect 100 436 104 444
rect 113 436 119 444
rect 100 433 119 436
rect 146 444 157 448
rect 146 437 148 444
rect 156 437 157 444
rect 146 433 157 437
rect 164 442 186 448
rect 164 436 167 442
rect 175 436 186 442
rect 164 433 186 436
rect 282 446 296 448
rect 282 440 285 446
rect 292 440 296 446
rect 282 433 296 440
rect 303 444 322 448
rect 303 436 307 444
rect 316 436 322 444
rect 303 433 322 436
rect 349 444 360 448
rect 349 437 351 444
rect 359 437 360 444
rect 349 433 360 437
rect 367 442 389 448
rect 367 436 370 442
rect 378 436 389 442
rect 367 433 389 436
rect 469 446 483 448
rect 469 440 472 446
rect 479 440 483 446
rect 469 433 483 440
rect 490 444 509 448
rect 490 436 494 444
rect 503 436 509 444
rect 490 433 509 436
rect 536 444 547 448
rect 536 437 538 444
rect 546 437 547 444
rect 536 433 547 437
rect 554 442 576 448
rect 554 436 557 442
rect 565 436 576 442
rect 554 433 576 436
rect 650 446 664 448
rect 650 440 653 446
rect 660 440 664 446
rect 650 433 664 440
rect 671 444 690 448
rect 671 436 675 444
rect 684 436 690 444
rect 671 433 690 436
rect 717 444 728 448
rect 717 437 719 444
rect 727 437 728 444
rect 717 433 728 437
rect 735 442 757 448
rect 735 436 738 442
rect 746 436 757 442
rect 735 433 757 436
rect 77 155 91 157
rect 77 149 80 155
rect 87 149 91 155
rect 77 142 91 149
rect 98 153 117 157
rect 98 145 102 153
rect 111 145 117 153
rect 98 142 117 145
rect 144 153 155 157
rect 144 146 146 153
rect 154 146 155 153
rect 144 142 155 146
rect 162 151 184 157
rect 162 145 165 151
rect 173 145 184 151
rect 162 142 184 145
rect 280 155 294 157
rect 280 149 283 155
rect 290 149 294 155
rect 280 142 294 149
rect 301 153 320 157
rect 301 145 305 153
rect 314 145 320 153
rect 301 142 320 145
rect 347 153 358 157
rect 347 146 349 153
rect 357 146 358 153
rect 347 142 358 146
rect 365 151 387 157
rect 365 145 368 151
rect 376 145 387 151
rect 365 142 387 145
rect 467 155 481 157
rect 467 149 470 155
rect 477 149 481 155
rect 467 142 481 149
rect 488 153 507 157
rect 488 145 492 153
rect 501 145 507 153
rect 488 142 507 145
rect 534 153 545 157
rect 534 146 536 153
rect 544 146 545 153
rect 534 142 545 146
rect 552 151 574 157
rect 552 145 555 151
rect 563 145 574 151
rect 552 142 574 145
rect 648 155 662 157
rect 648 149 651 155
rect 658 149 662 155
rect 648 142 662 149
rect 669 153 688 157
rect 669 145 673 153
rect 682 145 688 153
rect 669 142 688 145
rect 715 153 726 157
rect 715 146 717 153
rect 725 146 726 153
rect 715 142 726 146
rect 733 151 755 157
rect 733 145 736 151
rect 744 145 755 151
rect 733 142 755 145
rect 1990 214 2004 216
rect 1990 208 1993 214
rect 2000 208 2004 214
rect 1990 201 2004 208
rect 2011 212 2030 216
rect 2011 204 2015 212
rect 2024 204 2030 212
rect 2011 201 2030 204
rect 2057 212 2068 216
rect 2057 205 2059 212
rect 2067 205 2068 212
rect 2057 201 2068 205
rect 2075 210 2097 216
rect 2075 204 2078 210
rect 2086 204 2097 210
rect 2075 201 2097 204
rect 2127 215 2141 217
rect 2127 209 2130 215
rect 2137 209 2141 215
rect 2127 202 2141 209
rect 2148 213 2167 217
rect 2148 205 2152 213
rect 2161 205 2167 213
rect 2148 202 2167 205
rect 2194 213 2205 217
rect 2194 206 2196 213
rect 2204 206 2205 213
rect 2194 202 2205 206
rect 2212 211 2234 217
rect 2212 205 2215 211
rect 2223 205 2234 211
rect 2212 202 2234 205
rect 2298 197 2300 206
rect 2306 197 2308 206
rect 2317 197 2321 206
<< ndcontact >>
rect 55 1006 63 1013
rect 77 1003 87 1012
rect 118 1006 126 1014
rect 141 1005 149 1013
rect 258 1006 266 1013
rect 280 1003 290 1012
rect 321 1006 329 1014
rect 344 1005 352 1013
rect 445 1006 453 1013
rect 467 1003 477 1012
rect 508 1006 516 1014
rect 531 1005 539 1013
rect 626 1006 634 1013
rect 648 1003 658 1012
rect 689 1006 697 1014
rect 712 1005 720 1013
rect 61 671 69 678
rect 83 668 93 677
rect 124 671 132 679
rect 147 670 155 678
rect 264 671 272 678
rect 286 668 296 677
rect 327 671 335 679
rect 350 670 358 678
rect 451 671 459 678
rect 473 668 483 677
rect 514 671 522 679
rect 537 670 545 678
rect 632 671 640 678
rect 654 668 664 677
rect 695 671 703 679
rect 718 670 726 678
rect 1004 386 1012 393
rect 1026 383 1036 392
rect 1067 386 1075 394
rect 1090 385 1098 393
rect 1143 386 1151 394
rect 1163 384 1173 393
rect 1204 387 1212 395
rect 1227 386 1235 394
rect 81 354 89 361
rect 103 351 113 360
rect 144 354 152 362
rect 167 353 175 361
rect 284 354 292 361
rect 306 351 316 360
rect 347 354 355 362
rect 370 353 378 361
rect 471 354 479 361
rect 493 351 503 360
rect 534 354 542 362
rect 557 353 565 361
rect 652 354 660 361
rect 674 351 684 360
rect 715 354 723 362
rect 738 353 746 361
rect 2290 146 2298 155
rect 2308 146 2316 155
rect 1992 122 2000 129
rect 2014 119 2024 128
rect 2055 122 2063 130
rect 2078 121 2086 129
rect 2131 122 2139 130
rect 2151 120 2161 129
rect 2192 123 2200 131
rect 2215 122 2223 130
rect 79 63 87 70
rect 101 60 111 69
rect 142 63 150 71
rect 165 62 173 70
rect 282 63 290 70
rect 304 60 314 69
rect 345 63 353 71
rect 368 62 376 70
rect 469 63 477 70
rect 491 60 501 69
rect 532 63 540 71
rect 555 62 563 70
rect 650 63 658 70
rect 672 60 682 69
rect 713 63 721 71
rect 736 62 744 70
<< pdcontact >>
rect 56 1092 63 1098
rect 78 1088 87 1096
rect 122 1089 130 1096
rect 141 1088 149 1094
rect 259 1092 266 1098
rect 281 1088 290 1096
rect 325 1089 333 1096
rect 344 1088 352 1094
rect 446 1092 453 1098
rect 468 1088 477 1096
rect 512 1089 520 1096
rect 531 1088 539 1094
rect 627 1092 634 1098
rect 649 1088 658 1096
rect 693 1089 701 1096
rect 712 1088 720 1094
rect 62 757 69 763
rect 84 753 93 761
rect 128 754 136 761
rect 147 753 155 759
rect 265 757 272 763
rect 287 753 296 761
rect 331 754 339 761
rect 350 753 358 759
rect 452 757 459 763
rect 474 753 483 761
rect 518 754 526 761
rect 537 753 545 759
rect 633 757 640 763
rect 655 753 664 761
rect 699 754 707 761
rect 718 753 726 759
rect 1005 472 1012 478
rect 1027 468 1036 476
rect 1071 469 1079 476
rect 1090 468 1098 474
rect 1142 473 1149 479
rect 1164 469 1173 477
rect 1208 470 1216 477
rect 1227 469 1235 475
rect 82 440 89 446
rect 104 436 113 444
rect 148 437 156 444
rect 167 436 175 442
rect 285 440 292 446
rect 307 436 316 444
rect 351 437 359 444
rect 370 436 378 442
rect 472 440 479 446
rect 494 436 503 444
rect 538 437 546 444
rect 557 436 565 442
rect 653 440 660 446
rect 675 436 684 444
rect 719 437 727 444
rect 738 436 746 442
rect 80 149 87 155
rect 102 145 111 153
rect 146 146 154 153
rect 165 145 173 151
rect 283 149 290 155
rect 305 145 314 153
rect 349 146 357 153
rect 368 145 376 151
rect 470 149 477 155
rect 492 145 501 153
rect 536 146 544 153
rect 555 145 563 151
rect 651 149 658 155
rect 673 145 682 153
rect 717 146 725 153
rect 736 145 744 151
rect 1993 208 2000 214
rect 2015 204 2024 212
rect 2059 205 2067 212
rect 2078 204 2086 210
rect 2130 209 2137 215
rect 2152 205 2161 213
rect 2196 206 2204 213
rect 2215 205 2223 211
rect 2290 197 2298 206
rect 2308 197 2317 206
<< polysilicon >>
rect 4 1157 478 1165
rect 4 1154 138 1157
rect 0 1126 28 1137
rect 18 1050 28 1126
rect 67 1100 74 1103
rect 131 1100 138 1154
rect 270 1100 277 1103
rect 334 1100 341 1103
rect 457 1100 464 1157
rect 521 1100 528 1103
rect 638 1100 645 1133
rect 702 1100 709 1103
rect 67 1050 74 1085
rect 18 1042 74 1050
rect 18 1041 28 1042
rect 67 1015 74 1042
rect 131 1015 138 1085
rect 270 1015 277 1085
rect 334 1015 341 1085
rect 457 1015 464 1085
rect 521 1015 528 1085
rect 638 1015 645 1085
rect 702 1015 709 1085
rect 1114 1058 1120 1077
rect 67 956 74 1000
rect 131 995 138 1000
rect 270 956 277 1000
rect 334 971 341 1000
rect 457 996 464 1000
rect 521 972 528 1000
rect 638 996 645 1000
rect 67 949 277 956
rect 702 953 709 1000
rect 10 822 484 830
rect 10 819 144 822
rect 6 791 34 802
rect 24 715 34 791
rect 73 765 80 768
rect 137 765 144 819
rect 276 765 283 768
rect 340 765 347 768
rect 463 765 470 822
rect 527 765 534 768
rect 644 765 651 798
rect 708 765 715 768
rect 73 715 80 750
rect 24 707 80 715
rect 24 706 34 707
rect 73 680 80 707
rect 137 680 144 750
rect 276 680 283 750
rect 340 680 347 750
rect 463 680 470 750
rect 527 680 534 750
rect 644 680 651 750
rect 708 680 715 750
rect 73 621 80 665
rect 137 660 144 665
rect 276 621 283 665
rect 340 636 347 665
rect 463 661 470 665
rect 527 637 534 665
rect 644 661 651 665
rect 73 614 283 621
rect 708 618 715 665
rect 1114 553 1120 1049
rect 30 505 504 513
rect 30 502 164 505
rect 26 474 54 485
rect 44 398 54 474
rect 93 448 100 451
rect 157 448 164 502
rect 296 448 303 451
rect 360 448 367 451
rect 483 448 490 505
rect 547 448 554 451
rect 664 448 671 481
rect 1016 480 1023 483
rect 1080 480 1087 483
rect 1153 481 1160 484
rect 1217 481 1224 484
rect 728 448 735 451
rect 93 398 100 433
rect 44 390 100 398
rect 44 389 54 390
rect 93 363 100 390
rect 157 363 164 433
rect 296 363 303 433
rect 360 363 367 433
rect 483 363 490 433
rect 547 363 554 433
rect 664 363 671 433
rect 728 363 735 433
rect 1016 395 1023 465
rect 1080 395 1087 465
rect 1153 396 1160 466
rect 1217 396 1224 466
rect 1016 376 1023 380
rect 1080 375 1087 380
rect 1153 377 1160 381
rect 1217 376 1224 381
rect 93 304 100 348
rect 157 343 164 348
rect 296 304 303 348
rect 360 319 367 348
rect 483 344 490 348
rect 547 320 554 348
rect 664 344 671 348
rect 93 297 303 304
rect 728 301 735 348
rect 28 214 502 222
rect 28 211 162 214
rect 24 183 52 194
rect 42 107 52 183
rect 91 157 98 160
rect 155 157 162 211
rect 294 157 301 160
rect 358 157 365 160
rect 481 157 488 214
rect 545 157 552 160
rect 662 157 669 190
rect 726 157 733 160
rect 91 107 98 142
rect 42 99 98 107
rect 42 98 52 99
rect 91 72 98 99
rect 155 72 162 142
rect 294 72 301 142
rect 358 72 365 142
rect 481 72 488 142
rect 545 72 552 142
rect 662 72 669 142
rect 726 72 733 142
rect 1071 111 1077 349
rect 2004 216 2011 219
rect 2068 216 2075 219
rect 2141 217 2148 220
rect 2205 217 2212 220
rect 2300 206 2306 209
rect 2004 131 2011 201
rect 2068 131 2075 201
rect 2141 132 2148 202
rect 2205 132 2212 202
rect 2300 170 2306 197
rect 2305 163 2306 170
rect 2300 155 2306 163
rect 2300 143 2306 146
rect 2004 112 2011 116
rect 2068 111 2075 116
rect 2141 113 2148 117
rect 2205 112 2212 117
rect 1071 79 1077 104
rect 91 13 98 57
rect 155 52 162 57
rect 294 13 301 57
rect 358 28 365 57
rect 481 53 488 57
rect 545 29 552 57
rect 662 53 669 57
rect 91 6 301 13
rect 726 10 733 57
<< polycontact >>
rect 638 1133 645 1140
rect 1113 1049 1121 1058
rect 334 963 341 971
rect 521 964 528 972
rect 702 946 709 953
rect 644 798 651 805
rect 340 628 347 636
rect 527 629 534 637
rect 708 611 715 618
rect 664 481 671 488
rect 360 311 367 319
rect 547 312 554 320
rect 728 294 735 301
rect 662 190 669 197
rect 2300 163 2305 170
rect 1070 104 1078 111
rect 358 20 365 28
rect 545 21 552 29
rect 726 3 733 10
<< metal1 >>
rect 387 1140 646 1142
rect 73 1129 372 1139
rect 387 1133 638 1140
rect 645 1133 646 1140
rect 387 1132 646 1133
rect 122 1118 130 1129
rect 325 1118 333 1129
rect 56 1112 130 1118
rect 56 1098 63 1112
rect 122 1096 130 1112
rect 259 1112 333 1118
rect 259 1098 266 1112
rect 78 1057 87 1088
rect 325 1096 333 1112
rect 141 1067 149 1088
rect 140 1057 149 1067
rect 78 1054 149 1057
rect 281 1057 290 1088
rect 344 1057 352 1088
rect 281 1056 352 1057
rect 388 1056 397 1132
rect 512 1118 520 1127
rect 693 1118 701 1127
rect 446 1112 520 1118
rect 446 1098 453 1112
rect 512 1096 520 1112
rect 78 1049 175 1054
rect 281 1049 397 1056
rect 627 1112 701 1118
rect 627 1098 634 1112
rect 468 1057 477 1088
rect 693 1096 701 1112
rect 531 1057 539 1088
rect 468 1056 539 1057
rect 649 1057 658 1088
rect 712 1057 720 1088
rect 649 1056 720 1057
rect 726 1056 1113 1058
rect 468 1049 585 1056
rect 649 1049 1113 1056
rect 141 1045 175 1049
rect 77 1021 126 1029
rect 55 984 63 1006
rect 77 1012 87 1021
rect 118 1014 126 1021
rect 141 1013 149 1045
rect 164 972 175 1045
rect 344 1047 397 1049
rect 531 1047 585 1049
rect 280 1021 329 1029
rect 258 984 266 1006
rect 280 1012 290 1021
rect 321 1014 329 1021
rect 344 1013 352 1047
rect 467 1021 516 1029
rect 445 984 453 1006
rect 467 1012 477 1021
rect 508 1014 516 1021
rect 531 1013 539 1047
rect 164 971 521 972
rect 164 963 334 971
rect 341 964 521 971
rect 528 964 562 972
rect 341 963 562 964
rect 164 961 562 963
rect 573 953 585 1047
rect 712 1047 740 1049
rect 648 1021 697 1029
rect 626 984 634 1006
rect 648 1012 658 1021
rect 689 1014 697 1021
rect 712 1013 720 1047
rect 573 946 702 953
rect 709 946 742 953
rect 573 943 742 946
rect 393 805 652 807
rect 79 794 378 804
rect 393 798 644 805
rect 651 798 652 805
rect 393 797 652 798
rect 128 783 136 794
rect 331 783 339 794
rect 62 777 136 783
rect 62 763 69 777
rect 128 761 136 777
rect 265 777 339 783
rect 265 763 272 777
rect 84 722 93 753
rect 331 761 339 777
rect 147 732 155 753
rect 146 722 155 732
rect 84 719 155 722
rect 287 722 296 753
rect 350 722 358 753
rect 287 721 358 722
rect 394 721 403 797
rect 518 783 526 792
rect 699 783 707 792
rect 452 777 526 783
rect 452 763 459 777
rect 518 761 526 777
rect 84 714 181 719
rect 287 714 403 721
rect 633 777 707 783
rect 633 763 640 777
rect 474 722 483 753
rect 699 761 707 777
rect 537 722 545 753
rect 474 721 545 722
rect 655 722 664 753
rect 718 722 726 753
rect 824 722 833 723
rect 655 721 726 722
rect 744 721 833 722
rect 474 714 591 721
rect 655 714 833 721
rect 147 710 181 714
rect 83 686 132 694
rect 61 649 69 671
rect 83 677 93 686
rect 124 679 132 686
rect 147 678 155 710
rect 170 637 181 710
rect 350 712 403 714
rect 537 712 591 714
rect 286 686 335 694
rect 264 649 272 671
rect 286 677 296 686
rect 327 679 335 686
rect 350 678 358 712
rect 473 686 522 694
rect 451 649 459 671
rect 473 677 483 686
rect 514 679 522 686
rect 537 678 545 712
rect 170 636 527 637
rect 170 628 340 636
rect 347 629 527 636
rect 534 629 568 637
rect 347 628 568 629
rect 170 626 568 628
rect 579 618 591 712
rect 718 712 833 714
rect 654 686 703 694
rect 632 649 640 671
rect 654 677 664 686
rect 695 679 703 686
rect 718 678 726 712
rect 744 711 833 712
rect 579 611 708 618
rect 715 611 748 618
rect 579 608 748 611
rect 824 497 833 711
rect 1071 499 1079 503
rect 1208 499 1216 504
rect 1071 498 1216 499
rect 413 488 672 490
rect 824 489 951 497
rect 1005 494 1216 498
rect 1005 492 1079 494
rect 99 477 398 487
rect 413 481 664 488
rect 671 481 672 488
rect 413 480 672 481
rect 148 466 156 477
rect 351 466 359 477
rect 82 460 156 466
rect 82 446 89 460
rect 148 444 156 460
rect 285 460 359 466
rect 285 446 292 460
rect 104 405 113 436
rect 351 444 359 460
rect 167 415 175 436
rect 166 405 175 415
rect 104 402 175 405
rect 307 405 316 436
rect 370 405 378 436
rect 307 404 378 405
rect 414 404 423 480
rect 1005 478 1012 492
rect 538 466 546 475
rect 719 466 727 475
rect 1071 476 1079 492
rect 472 460 546 466
rect 472 446 479 460
rect 538 444 546 460
rect 104 397 201 402
rect 307 397 423 404
rect 653 460 727 466
rect 653 446 660 460
rect 494 405 503 436
rect 719 444 727 460
rect 557 405 565 436
rect 494 404 565 405
rect 1142 493 1216 494
rect 1142 479 1149 493
rect 675 405 684 436
rect 738 405 746 436
rect 1027 437 1036 468
rect 1208 477 1216 493
rect 1090 437 1098 468
rect 1027 435 1098 437
rect 1164 438 1173 469
rect 1227 438 1235 469
rect 1164 436 1235 438
rect 1164 435 1236 436
rect 1027 434 1099 435
rect 1109 434 1248 435
rect 1027 430 1248 434
rect 1027 429 1173 430
rect 1090 428 1173 429
rect 1090 426 1111 428
rect 1227 426 1248 430
rect 675 404 746 405
rect 494 397 611 404
rect 675 397 951 404
rect 167 393 201 397
rect 103 369 152 377
rect 81 332 89 354
rect 103 360 113 369
rect 144 362 152 369
rect 167 361 175 393
rect 190 320 201 393
rect 370 395 423 397
rect 557 395 611 397
rect 306 369 355 377
rect 284 332 292 354
rect 306 360 316 369
rect 347 362 355 369
rect 370 361 378 395
rect 493 369 542 377
rect 471 332 479 354
rect 493 360 503 369
rect 534 362 542 369
rect 557 361 565 395
rect 190 319 547 320
rect 190 311 360 319
rect 367 312 547 319
rect 554 312 588 320
rect 367 311 588 312
rect 190 309 588 311
rect 599 301 611 395
rect 738 395 951 397
rect 674 369 723 377
rect 652 332 660 354
rect 674 360 684 369
rect 715 362 723 369
rect 738 361 746 395
rect 755 394 951 395
rect 1026 401 1075 409
rect 1004 364 1012 386
rect 1026 392 1036 401
rect 1067 394 1075 401
rect 1090 403 1151 412
rect 1090 393 1098 403
rect 1143 394 1151 403
rect 1163 402 1212 410
rect 1163 393 1173 402
rect 1204 395 1212 402
rect 1227 394 1235 426
rect 599 294 728 301
rect 735 294 768 301
rect 599 291 768 294
rect 2059 235 2067 239
rect 2196 235 2204 240
rect 2059 234 2204 235
rect 1993 230 2204 234
rect 1993 228 2067 230
rect 1993 214 2000 228
rect 2059 212 2067 228
rect 2130 229 2204 230
rect 2130 215 2137 229
rect 411 197 670 199
rect 97 186 396 196
rect 411 190 662 197
rect 669 190 670 197
rect 411 189 670 190
rect 146 175 154 186
rect 349 175 357 186
rect 80 169 154 175
rect 80 155 87 169
rect 146 153 154 169
rect 283 169 357 175
rect 283 155 290 169
rect 102 114 111 145
rect 349 153 357 169
rect 165 124 173 145
rect 164 114 173 124
rect 102 111 173 114
rect 305 114 314 145
rect 368 114 376 145
rect 305 113 376 114
rect 412 113 421 189
rect 536 175 544 184
rect 717 175 725 184
rect 470 169 544 175
rect 470 155 477 169
rect 536 153 544 169
rect 102 106 199 111
rect 305 106 421 113
rect 651 169 725 175
rect 651 155 658 169
rect 492 114 501 145
rect 717 153 725 169
rect 2015 173 2024 204
rect 2196 213 2204 229
rect 2078 173 2086 204
rect 2015 171 2086 173
rect 2152 174 2161 205
rect 2291 206 2298 222
rect 2215 174 2223 205
rect 2152 172 2223 174
rect 2152 171 2224 172
rect 2015 170 2087 171
rect 2097 170 2236 171
rect 2015 166 2300 170
rect 2015 165 2161 166
rect 2078 164 2161 165
rect 2078 162 2099 164
rect 2215 163 2300 166
rect 2215 162 2236 163
rect 555 114 563 145
rect 492 113 563 114
rect 673 114 682 145
rect 736 114 744 145
rect 2014 137 2063 145
rect 673 113 744 114
rect 492 106 609 113
rect 673 112 764 113
rect 673 111 1078 112
rect 673 106 1070 111
rect 165 102 199 106
rect 101 78 150 86
rect 79 41 87 63
rect 101 69 111 78
rect 142 71 150 78
rect 165 70 173 102
rect 188 29 199 102
rect 368 104 421 106
rect 555 104 609 106
rect 304 78 353 86
rect 282 41 290 63
rect 304 69 314 78
rect 345 71 353 78
rect 368 70 376 104
rect 491 78 540 86
rect 469 41 477 63
rect 491 69 501 78
rect 532 71 540 78
rect 555 70 563 104
rect 188 28 545 29
rect 188 20 358 28
rect 365 21 545 28
rect 552 21 586 29
rect 365 20 586 21
rect 188 18 586 20
rect 597 10 609 104
rect 736 104 1070 106
rect 672 78 721 86
rect 650 41 658 63
rect 672 69 682 78
rect 713 71 721 78
rect 736 70 744 104
rect 1992 100 2000 122
rect 2014 128 2024 137
rect 2055 130 2063 137
rect 2078 139 2139 148
rect 2078 129 2086 139
rect 2131 130 2139 139
rect 2151 138 2200 146
rect 2151 129 2161 138
rect 2192 131 2200 138
rect 2215 130 2223 162
rect 2308 155 2316 197
rect 2291 136 2298 146
rect 597 3 726 10
rect 733 3 766 10
rect 597 0 766 3
<< labels >>
rlabel metal1 2031 229 2032 233 5 vdd
rlabel metal1 1998 104 1999 108 1 gnd
rlabel metal1 2168 230 2169 234 5 vdd
rlabel metal1 1180 494 1181 498 5 vdd
rlabel metal1 1010 368 1011 372 1 gnd
rlabel metal1 1043 493 1044 497 5 vdd
rlabel metal1 689 170 690 174 5 vdd
rlabel metal1 656 45 657 49 1 gnd
rlabel metal1 508 170 509 174 5 vdd
rlabel metal1 475 45 476 49 1 gnd
rlabel metal1 321 170 322 174 5 vdd
rlabel metal1 288 45 289 49 1 gnd
rlabel metal1 118 170 119 174 5 vdd
rlabel metal1 85 45 86 49 1 gnd
rlabel metal1 691 461 692 465 5 vdd
rlabel metal1 658 336 659 340 1 gnd
rlabel metal1 510 461 511 465 5 vdd
rlabel metal1 477 336 478 340 1 gnd
rlabel metal1 323 461 324 465 5 vdd
rlabel metal1 290 336 291 340 1 gnd
rlabel metal1 120 461 121 465 5 vdd
rlabel metal1 87 336 88 340 1 gnd
rlabel metal1 671 778 672 782 5 vdd
rlabel metal1 638 653 639 657 1 gnd
rlabel metal1 490 778 491 782 5 vdd
rlabel metal1 457 653 458 657 1 gnd
rlabel metal1 303 778 304 782 5 vdd
rlabel metal1 270 653 271 657 1 gnd
rlabel metal1 100 778 101 782 5 vdd
rlabel metal1 67 653 68 657 1 gnd
rlabel metal1 665 1113 666 1117 5 vdd
rlabel metal1 632 988 633 992 1 gnd
rlabel metal1 484 1113 485 1117 5 vdd
rlabel metal1 451 988 452 992 1 gnd
rlabel metal1 297 1113 298 1117 5 vdd
rlabel metal1 264 988 265 992 1 gnd
rlabel metal1 94 1113 95 1117 5 vdd
rlabel metal1 61 988 62 992 1 gnd
rlabel metal1 2292 215 2295 218 1 vdd
rlabel metal1 2292 138 2296 140 1 gnd
<< end >>
