magic
tech scmos
timestamp 1700463188
<< nwell >>
rect 0 96 131 137
rect 169 85 235 127
rect 2 -102 133 -61
rect 171 -113 237 -71
rect 2 -300 133 -259
rect 171 -311 237 -269
rect 2 -495 133 -454
rect 171 -506 237 -464
<< ntransistor >>
rect 26 26 33 41
rect 90 26 97 41
rect 199 20 207 36
rect 28 -172 35 -157
rect 92 -172 99 -157
rect 201 -178 209 -162
rect 28 -370 35 -355
rect 92 -370 99 -355
rect 201 -376 209 -360
rect 28 -565 35 -550
rect 92 -565 99 -550
rect 201 -571 209 -555
<< ptransistor >>
rect 26 111 33 126
rect 90 111 97 126
rect 199 98 207 114
rect 28 -87 35 -72
rect 92 -87 99 -72
rect 201 -100 209 -84
rect 28 -285 35 -270
rect 92 -285 99 -270
rect 201 -298 209 -282
rect 28 -480 35 -465
rect 92 -480 99 -465
rect 201 -493 209 -477
<< ndiffusion >>
rect 12 39 26 41
rect 12 32 14 39
rect 22 32 26 39
rect 12 26 26 32
rect 33 38 52 41
rect 33 29 36 38
rect 46 29 52 38
rect 33 26 52 29
rect 71 40 90 41
rect 71 32 77 40
rect 85 32 90 40
rect 71 26 90 32
rect 97 39 111 41
rect 97 31 100 39
rect 108 31 111 39
rect 97 26 111 31
rect 182 32 199 36
rect 182 22 184 32
rect 194 22 199 32
rect 182 20 199 22
rect 207 33 222 36
rect 207 23 209 33
rect 219 23 222 33
rect 207 20 222 23
rect 14 -159 28 -157
rect 14 -166 16 -159
rect 24 -166 28 -159
rect 14 -172 28 -166
rect 35 -160 54 -157
rect 35 -169 38 -160
rect 48 -169 54 -160
rect 35 -172 54 -169
rect 73 -158 92 -157
rect 73 -166 79 -158
rect 87 -166 92 -158
rect 73 -172 92 -166
rect 99 -159 113 -157
rect 99 -167 102 -159
rect 110 -167 113 -159
rect 99 -172 113 -167
rect 184 -166 201 -162
rect 184 -176 186 -166
rect 196 -176 201 -166
rect 184 -178 201 -176
rect 209 -165 224 -162
rect 209 -175 211 -165
rect 221 -175 224 -165
rect 209 -178 224 -175
rect 14 -357 28 -355
rect 14 -364 16 -357
rect 24 -364 28 -357
rect 14 -370 28 -364
rect 35 -358 54 -355
rect 35 -367 38 -358
rect 48 -367 54 -358
rect 35 -370 54 -367
rect 73 -356 92 -355
rect 73 -364 79 -356
rect 87 -364 92 -356
rect 73 -370 92 -364
rect 99 -357 113 -355
rect 99 -365 102 -357
rect 110 -365 113 -357
rect 99 -370 113 -365
rect 184 -364 201 -360
rect 184 -374 186 -364
rect 196 -374 201 -364
rect 184 -376 201 -374
rect 209 -363 224 -360
rect 209 -373 211 -363
rect 221 -373 224 -363
rect 209 -376 224 -373
rect 14 -552 28 -550
rect 14 -559 16 -552
rect 24 -559 28 -552
rect 14 -565 28 -559
rect 35 -553 54 -550
rect 35 -562 38 -553
rect 48 -562 54 -553
rect 35 -565 54 -562
rect 73 -551 92 -550
rect 73 -559 79 -551
rect 87 -559 92 -551
rect 73 -565 92 -559
rect 99 -552 113 -550
rect 99 -560 102 -552
rect 110 -560 113 -552
rect 99 -565 113 -560
rect 184 -559 201 -555
rect 184 -569 186 -559
rect 196 -569 201 -559
rect 184 -571 201 -569
rect 209 -558 224 -555
rect 209 -568 211 -558
rect 221 -568 224 -558
rect 209 -571 224 -568
<< pdiffusion >>
rect 12 124 26 126
rect 12 118 15 124
rect 22 118 26 124
rect 12 111 26 118
rect 33 122 52 126
rect 33 114 37 122
rect 46 114 52 122
rect 33 111 52 114
rect 79 122 90 126
rect 79 115 81 122
rect 89 115 90 122
rect 79 111 90 115
rect 97 120 119 126
rect 97 114 100 120
rect 108 114 119 120
rect 97 111 119 114
rect 183 104 185 114
rect 195 104 199 114
rect 183 98 199 104
rect 207 111 223 114
rect 207 101 209 111
rect 219 101 223 111
rect 207 98 223 101
rect 14 -74 28 -72
rect 14 -80 17 -74
rect 24 -80 28 -74
rect 14 -87 28 -80
rect 35 -76 54 -72
rect 35 -84 39 -76
rect 48 -84 54 -76
rect 35 -87 54 -84
rect 81 -76 92 -72
rect 81 -83 83 -76
rect 91 -83 92 -76
rect 81 -87 92 -83
rect 99 -78 121 -72
rect 99 -84 102 -78
rect 110 -84 121 -78
rect 99 -87 121 -84
rect 185 -94 187 -84
rect 197 -94 201 -84
rect 185 -100 201 -94
rect 209 -87 225 -84
rect 209 -97 211 -87
rect 221 -97 225 -87
rect 209 -100 225 -97
rect 14 -272 28 -270
rect 14 -278 17 -272
rect 24 -278 28 -272
rect 14 -285 28 -278
rect 35 -274 54 -270
rect 35 -282 39 -274
rect 48 -282 54 -274
rect 35 -285 54 -282
rect 81 -274 92 -270
rect 81 -281 83 -274
rect 91 -281 92 -274
rect 81 -285 92 -281
rect 99 -276 121 -270
rect 99 -282 102 -276
rect 110 -282 121 -276
rect 99 -285 121 -282
rect 185 -292 187 -282
rect 197 -292 201 -282
rect 185 -298 201 -292
rect 209 -285 225 -282
rect 209 -295 211 -285
rect 221 -295 225 -285
rect 209 -298 225 -295
rect 14 -467 28 -465
rect 14 -473 17 -467
rect 24 -473 28 -467
rect 14 -480 28 -473
rect 35 -469 54 -465
rect 35 -477 39 -469
rect 48 -477 54 -469
rect 35 -480 54 -477
rect 81 -469 92 -465
rect 81 -476 83 -469
rect 91 -476 92 -469
rect 81 -480 92 -476
rect 99 -471 121 -465
rect 99 -477 102 -471
rect 110 -477 121 -471
rect 99 -480 121 -477
rect 185 -487 187 -477
rect 197 -487 201 -477
rect 185 -493 201 -487
rect 209 -480 225 -477
rect 209 -490 211 -480
rect 221 -490 225 -480
rect 209 -493 225 -490
<< ndcontact >>
rect 14 32 22 39
rect 36 29 46 38
rect 77 32 85 40
rect 100 31 108 39
rect 184 22 194 32
rect 209 23 219 33
rect 16 -166 24 -159
rect 38 -169 48 -160
rect 79 -166 87 -158
rect 102 -167 110 -159
rect 186 -176 196 -166
rect 211 -175 221 -165
rect 16 -364 24 -357
rect 38 -367 48 -358
rect 79 -364 87 -356
rect 102 -365 110 -357
rect 186 -374 196 -364
rect 211 -373 221 -363
rect 16 -559 24 -552
rect 38 -562 48 -553
rect 79 -559 87 -551
rect 102 -560 110 -552
rect 186 -569 196 -559
rect 211 -568 221 -558
<< pdcontact >>
rect 15 118 22 124
rect 37 114 46 122
rect 81 115 89 122
rect 100 114 108 120
rect 185 104 195 114
rect 209 101 219 111
rect 17 -80 24 -74
rect 39 -84 48 -76
rect 83 -83 91 -76
rect 102 -84 110 -78
rect 187 -94 197 -84
rect 211 -97 221 -87
rect 17 -278 24 -272
rect 39 -282 48 -274
rect 83 -281 91 -274
rect 102 -282 110 -276
rect 187 -292 197 -282
rect 211 -295 221 -285
rect 17 -473 24 -467
rect 39 -477 48 -469
rect 83 -476 91 -469
rect 102 -477 110 -471
rect 187 -487 197 -477
rect 211 -490 221 -480
<< polysilicon >>
rect -344 159 97 167
rect -344 158 -56 159
rect -344 3 -327 158
rect 26 126 33 129
rect 90 126 97 159
rect 199 114 207 120
rect 26 41 33 111
rect 90 41 97 111
rect 199 67 207 98
rect 165 66 207 67
rect 175 57 207 66
rect 199 36 207 57
rect -281 -4 -71 -3
rect 26 -4 33 26
rect 90 21 97 26
rect 199 12 207 20
rect -281 -12 34 -4
rect -281 -22 -266 -12
rect -211 -31 97 -30
rect -197 -39 99 -31
rect 28 -72 35 -69
rect 92 -72 99 -39
rect 201 -84 209 -78
rect 28 -157 35 -87
rect 92 -157 99 -87
rect 201 -131 209 -100
rect 167 -132 209 -131
rect 177 -141 209 -132
rect 201 -162 209 -141
rect -194 -202 -63 -201
rect 28 -202 35 -172
rect 92 -177 99 -172
rect 201 -186 209 -178
rect -194 -210 36 -202
rect -341 -237 99 -229
rect -340 -324 -326 -237
rect 28 -270 35 -267
rect 92 -270 99 -237
rect 201 -282 209 -276
rect -327 -338 -326 -324
rect 28 -355 35 -285
rect 92 -355 99 -285
rect 201 -329 209 -298
rect 167 -330 209 -329
rect 177 -339 209 -330
rect 201 -360 209 -339
rect -150 -404 -149 -390
rect 28 -400 35 -370
rect 92 -375 99 -370
rect 201 -384 209 -376
rect -161 -423 -149 -404
rect -66 -408 36 -400
rect -161 -424 -50 -423
rect -161 -432 99 -424
rect 28 -465 35 -462
rect 92 -465 99 -432
rect 201 -477 209 -471
rect 28 -550 35 -480
rect 92 -550 99 -480
rect 201 -524 209 -493
rect 167 -525 209 -524
rect 177 -534 209 -525
rect 201 -555 209 -534
rect 28 -595 35 -565
rect 92 -570 99 -565
rect 201 -579 209 -571
rect -79 -603 -78 -595
rect -59 -603 36 -595
<< polycontact >>
rect 164 56 175 66
rect -344 -11 -325 3
rect -282 -38 -266 -22
rect -211 -40 -197 -31
rect 166 -142 177 -132
rect -208 -210 -194 -201
rect -341 -339 -327 -324
rect 166 -340 177 -330
rect -161 -404 -150 -390
rect -79 -408 -66 -400
rect 166 -535 177 -525
rect -78 -604 -59 -595
<< metal1 >>
rect 81 144 89 149
rect 15 138 89 144
rect 15 124 22 138
rect 81 122 89 138
rect 221 134 229 142
rect 186 128 229 134
rect 37 83 46 114
rect 186 114 194 128
rect 100 83 108 114
rect 37 81 108 83
rect 37 80 109 81
rect 37 75 134 80
rect 100 71 134 75
rect 36 47 85 55
rect 14 10 22 32
rect 36 38 46 47
rect 77 40 85 47
rect 100 39 108 71
rect 123 66 134 71
rect 209 68 219 101
rect 123 56 164 66
rect 209 59 243 68
rect 209 33 219 59
rect 185 6 194 22
rect -479 3 -327 4
rect -479 -10 -344 3
rect 185 0 220 6
rect -479 -37 -282 -23
rect -349 -38 -282 -37
rect -266 -38 -265 -23
rect -212 -40 -211 -31
rect -212 -48 -198 -40
rect -352 -49 -197 -48
rect -479 -63 -197 -49
rect 83 -54 91 -49
rect 17 -60 91 -54
rect 17 -74 24 -60
rect -479 -92 -194 -79
rect 83 -76 91 -60
rect 223 -64 231 -56
rect -479 -93 -327 -92
rect -208 -201 -194 -92
rect 188 -70 231 -64
rect 39 -115 48 -84
rect 188 -84 196 -70
rect 102 -115 110 -84
rect 39 -117 110 -115
rect 39 -118 111 -117
rect 39 -123 136 -118
rect 102 -127 136 -123
rect 38 -151 87 -143
rect 16 -188 24 -166
rect 38 -160 48 -151
rect 79 -158 87 -151
rect 102 -159 110 -127
rect 125 -132 136 -127
rect 211 -130 221 -97
rect 125 -142 166 -132
rect 211 -139 246 -130
rect 211 -165 221 -139
rect 187 -192 196 -176
rect 187 -198 222 -192
rect -208 -211 -194 -210
rect 83 -252 91 -247
rect 17 -258 91 -252
rect 17 -272 24 -258
rect 83 -274 91 -258
rect 223 -262 231 -254
rect 188 -268 231 -262
rect 39 -313 48 -282
rect 188 -282 196 -268
rect 102 -313 110 -282
rect 39 -315 110 -313
rect 39 -316 111 -315
rect 39 -321 136 -316
rect -479 -338 -341 -324
rect 102 -325 136 -321
rect 38 -349 87 -341
rect -479 -369 -66 -355
rect -479 -404 -161 -390
rect -336 -405 -150 -404
rect -79 -400 -66 -369
rect 16 -386 24 -364
rect 38 -358 48 -349
rect 79 -356 87 -349
rect 102 -357 110 -325
rect 125 -330 136 -325
rect 211 -328 221 -295
rect 125 -340 166 -330
rect 211 -337 248 -328
rect 211 -363 221 -337
rect 187 -390 196 -374
rect 187 -396 222 -390
rect -479 -439 -327 -425
rect -342 -594 -327 -439
rect 83 -447 91 -442
rect 17 -453 91 -447
rect 17 -467 24 -453
rect 83 -469 91 -453
rect 223 -457 231 -449
rect 188 -463 231 -457
rect 39 -508 48 -477
rect 188 -477 196 -463
rect 102 -508 110 -477
rect 39 -510 110 -508
rect 39 -511 111 -510
rect 39 -516 136 -511
rect 102 -520 136 -516
rect 38 -544 87 -536
rect 16 -581 24 -559
rect 38 -553 48 -544
rect 79 -551 87 -544
rect 102 -552 110 -520
rect 125 -525 136 -520
rect 211 -523 221 -490
rect 125 -535 166 -525
rect 211 -532 248 -523
rect 211 -558 221 -532
rect 187 -585 196 -569
rect 187 -591 222 -585
rect -342 -595 -59 -594
rect -342 -604 -78 -595
<< labels >>
rlabel metal1 204 131 206 133 5 vdd
rlabel metal1 214 2 216 4 1 gnd
rlabel metal1 53 139 54 143 5 vdd
rlabel metal1 20 14 21 18 1 gnd
rlabel metal1 206 -67 208 -65 5 vdd
rlabel metal1 216 -196 218 -194 1 gnd
rlabel metal1 55 -59 56 -55 5 vdd
rlabel metal1 22 -184 23 -180 1 gnd
rlabel metal1 206 -265 208 -263 5 vdd
rlabel metal1 216 -394 218 -392 1 gnd
rlabel metal1 55 -257 56 -253 5 vdd
rlabel metal1 22 -382 23 -378 1 gnd
rlabel metal1 206 -460 208 -458 5 vdd
rlabel metal1 216 -589 218 -587 1 gnd
rlabel metal1 55 -452 56 -448 5 vdd
rlabel metal1 22 -577 23 -573 1 gnd
rlabel metal1 -472 -4 -469 0 1 a0
rlabel metal1 -448 -34 -445 -30 1 b0
rlabel metal1 -400 -59 -397 -55 1 a1
rlabel metal1 -418 -88 -415 -84 1 b1
rlabel metal1 -435 -329 -432 -325 1 a2
rlabel metal1 -400 -368 -397 -364 1 b2
rlabel metal1 -449 -399 -446 -395 1 a3
rlabel metal1 -464 -434 -461 -430 1 b3
rlabel metal1 237 61 239 62 1 y0
rlabel metal1 230 -134 232 -133 1 y1
rlabel metal1 239 -334 241 -333 1 y2
rlabel metal1 236 -530 238 -529 1 y3
<< end >>
