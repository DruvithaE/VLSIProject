magic
tech scmos
timestamp 1700933555
<< nwell >>
rect 360 1973 491 2014
rect 529 1962 595 2004
rect 277 1899 324 1924
rect 1327 1896 1547 1921
rect 360 1844 491 1845
rect 360 1804 554 1844
rect 584 1807 650 1849
rect 491 1803 554 1804
rect 279 1737 326 1762
rect 340 1685 471 1686
rect 340 1684 529 1685
rect 340 1683 542 1684
rect 340 1645 597 1683
rect 604 1646 670 1688
rect 471 1644 597 1645
rect 535 1643 597 1644
rect 539 1642 597 1643
rect 278 1582 325 1607
rect 349 1466 480 1467
rect 349 1465 538 1466
rect 349 1464 551 1465
rect 349 1463 610 1464
rect 674 1463 740 1468
rect 349 1426 740 1463
rect 480 1425 676 1426
rect 544 1424 676 1425
rect 548 1423 676 1424
rect 607 1422 676 1423
rect 657 1421 676 1422
rect 278 1350 325 1375
rect 229 1036 360 1077
rect 432 1036 563 1077
rect 619 1036 750 1077
rect 800 1036 931 1077
rect 963 1032 1010 1057
rect 235 747 366 788
rect 438 747 569 788
rect 625 747 756 788
rect 806 747 937 788
rect 965 740 1012 765
rect 255 430 386 471
rect 458 430 589 471
rect 645 430 776 471
rect 826 430 957 471
rect 1178 462 1309 503
rect 1315 463 1446 504
rect 1452 459 1499 484
rect 990 423 1037 448
rect 253 139 384 180
rect 456 139 587 180
rect 643 139 774 180
rect 824 139 955 180
rect 999 132 1046 157
rect 306 -293 437 -252
rect 475 -304 541 -262
rect 223 -367 270 -342
rect 1387 -370 1607 -345
rect 306 -422 437 -421
rect 306 -462 500 -422
rect 530 -459 596 -417
rect 437 -463 500 -462
rect 225 -529 272 -504
rect 286 -581 417 -580
rect 286 -582 475 -581
rect 286 -583 488 -582
rect 286 -621 543 -583
rect 550 -620 616 -578
rect 417 -622 543 -621
rect 481 -623 543 -622
rect 485 -624 543 -623
rect 224 -684 271 -659
rect 295 -800 426 -799
rect 295 -801 484 -800
rect 295 -802 497 -801
rect 295 -803 556 -802
rect 620 -803 686 -798
rect 295 -840 686 -803
rect 426 -841 622 -840
rect 490 -842 622 -841
rect 494 -843 622 -842
rect 553 -844 622 -843
rect 603 -845 622 -844
rect 224 -916 271 -891
<< ntransistor >>
rect 386 1903 393 1918
rect 450 1903 457 1918
rect 559 1897 567 1913
rect 295 1856 301 1865
rect 1349 1842 1355 1853
rect 1390 1842 1396 1853
rect 1429 1842 1435 1853
rect 1472 1842 1478 1853
rect 1514 1842 1520 1853
rect 386 1734 393 1749
rect 450 1734 457 1749
rect 513 1733 520 1748
rect 614 1742 622 1758
rect 297 1694 303 1703
rect 366 1575 373 1590
rect 430 1575 437 1590
rect 493 1574 500 1589
rect 561 1572 568 1587
rect 634 1581 642 1597
rect 296 1539 302 1548
rect 375 1356 382 1371
rect 439 1356 446 1371
rect 502 1355 509 1370
rect 570 1353 577 1368
rect 629 1352 636 1367
rect 704 1361 712 1377
rect 296 1307 302 1316
rect 981 989 987 998
rect 255 966 262 981
rect 319 966 326 981
rect 458 966 465 981
rect 522 966 529 981
rect 645 966 652 981
rect 709 966 716 981
rect 826 966 833 981
rect 890 966 897 981
rect 983 697 989 706
rect 261 677 268 692
rect 325 677 332 692
rect 464 677 471 692
rect 528 677 535 692
rect 651 677 658 692
rect 715 677 722 692
rect 832 677 839 692
rect 896 677 903 692
rect 1008 380 1014 389
rect 281 360 288 375
rect 345 360 352 375
rect 484 360 491 375
rect 548 360 555 375
rect 671 360 678 375
rect 735 360 742 375
rect 852 360 859 375
rect 916 360 923 375
rect 1017 89 1023 98
rect 279 69 286 84
rect 343 69 350 84
rect 482 69 489 84
rect 546 69 553 84
rect 669 69 676 84
rect 733 69 740 84
rect 850 69 857 84
rect 914 69 921 84
rect 332 -363 339 -348
rect 396 -363 403 -348
rect 505 -369 513 -353
rect 241 -410 247 -401
rect 332 -532 339 -517
rect 396 -532 403 -517
rect 459 -533 466 -518
rect 560 -524 568 -508
rect 1470 416 1476 425
rect 1204 392 1211 407
rect 1268 392 1275 407
rect 1341 393 1348 408
rect 1405 393 1412 408
rect 243 -572 249 -563
rect 312 -691 319 -676
rect 376 -691 383 -676
rect 439 -692 446 -677
rect 507 -694 514 -679
rect 580 -685 588 -669
rect 242 -727 248 -718
rect 321 -910 328 -895
rect 385 -910 392 -895
rect 448 -911 455 -896
rect 516 -913 523 -898
rect 575 -914 582 -899
rect 650 -905 658 -889
rect 1409 -424 1415 -413
rect 1450 -424 1456 -413
rect 1489 -424 1495 -413
rect 1532 -424 1538 -413
rect 1574 -424 1580 -413
rect 242 -959 248 -950
<< ptransistor >>
rect 386 1988 393 2003
rect 450 1988 457 2003
rect 559 1975 567 1991
rect 295 1907 301 1916
rect 1349 1903 1355 1914
rect 1390 1903 1396 1914
rect 1429 1903 1435 1914
rect 1472 1903 1478 1914
rect 1514 1903 1520 1914
rect 386 1819 393 1834
rect 450 1819 457 1834
rect 297 1745 303 1754
rect 513 1818 520 1833
rect 614 1820 622 1836
rect 366 1660 373 1675
rect 430 1660 437 1675
rect 296 1590 302 1599
rect 493 1659 500 1674
rect 561 1657 568 1672
rect 634 1659 642 1675
rect 375 1441 382 1456
rect 439 1441 446 1456
rect 502 1440 509 1455
rect 296 1358 302 1367
rect 570 1438 577 1453
rect 629 1437 636 1452
rect 704 1439 712 1455
rect 255 1051 262 1066
rect 319 1051 326 1066
rect 458 1051 465 1066
rect 522 1051 529 1066
rect 645 1051 652 1066
rect 709 1051 716 1066
rect 826 1051 833 1066
rect 890 1051 897 1066
rect 981 1040 987 1049
rect 261 762 268 777
rect 325 762 332 777
rect 464 762 471 777
rect 528 762 535 777
rect 651 762 658 777
rect 715 762 722 777
rect 832 762 839 777
rect 896 762 903 777
rect 983 748 989 757
rect 281 445 288 460
rect 345 445 352 460
rect 484 445 491 460
rect 548 445 555 460
rect 671 445 678 460
rect 735 445 742 460
rect 852 445 859 460
rect 916 445 923 460
rect 1008 431 1014 440
rect 279 154 286 169
rect 343 154 350 169
rect 482 154 489 169
rect 546 154 553 169
rect 669 154 676 169
rect 733 154 740 169
rect 850 154 857 169
rect 914 154 921 169
rect 1017 140 1023 149
rect 332 -278 339 -263
rect 396 -278 403 -263
rect 505 -291 513 -275
rect 241 -359 247 -350
rect 332 -447 339 -432
rect 396 -447 403 -432
rect 243 -521 249 -512
rect 459 -448 466 -433
rect 560 -446 568 -430
rect 1204 477 1211 492
rect 1268 477 1275 492
rect 1341 478 1348 493
rect 1405 478 1412 493
rect 1470 467 1476 476
rect 312 -606 319 -591
rect 376 -606 383 -591
rect 242 -676 248 -667
rect 439 -607 446 -592
rect 507 -609 514 -594
rect 580 -607 588 -591
rect 321 -825 328 -810
rect 385 -825 392 -810
rect 448 -826 455 -811
rect 242 -908 248 -899
rect 516 -828 523 -813
rect 575 -829 582 -814
rect 650 -827 658 -811
rect 1409 -363 1415 -352
rect 1450 -363 1456 -352
rect 1489 -363 1495 -352
rect 1532 -363 1538 -352
rect 1574 -363 1580 -352
<< ndiffusion >>
rect 372 1916 386 1918
rect 372 1909 374 1916
rect 382 1909 386 1916
rect 372 1903 386 1909
rect 393 1915 412 1918
rect 393 1906 396 1915
rect 406 1906 412 1915
rect 393 1903 412 1906
rect 431 1917 450 1918
rect 431 1909 437 1917
rect 445 1909 450 1917
rect 431 1903 450 1909
rect 457 1916 471 1918
rect 457 1908 460 1916
rect 468 1908 471 1916
rect 457 1903 471 1908
rect 542 1909 559 1913
rect 542 1899 544 1909
rect 554 1899 559 1909
rect 542 1897 559 1899
rect 567 1910 582 1913
rect 567 1900 569 1910
rect 579 1900 582 1910
rect 567 1897 582 1900
rect 293 1856 295 1865
rect 301 1856 303 1865
rect 311 1856 316 1865
rect 1338 1850 1349 1853
rect 1338 1845 1340 1850
rect 1346 1845 1349 1850
rect 1338 1842 1349 1845
rect 1355 1851 1371 1853
rect 1355 1845 1359 1851
rect 1366 1845 1371 1851
rect 1355 1842 1371 1845
rect 1376 1850 1390 1853
rect 1376 1845 1380 1850
rect 1386 1845 1390 1850
rect 1376 1842 1390 1845
rect 1396 1851 1409 1853
rect 1396 1845 1399 1851
rect 1406 1845 1409 1851
rect 1396 1842 1409 1845
rect 1415 1850 1429 1853
rect 1415 1844 1419 1850
rect 1425 1844 1429 1850
rect 1415 1842 1429 1844
rect 1435 1852 1448 1853
rect 1435 1845 1438 1852
rect 1445 1845 1448 1852
rect 1435 1842 1448 1845
rect 1458 1850 1472 1853
rect 1458 1844 1462 1850
rect 1468 1844 1472 1850
rect 1458 1842 1472 1844
rect 1478 1851 1491 1853
rect 1478 1845 1480 1851
rect 1487 1845 1491 1851
rect 1478 1842 1491 1845
rect 1498 1850 1514 1853
rect 1498 1845 1504 1850
rect 1510 1845 1514 1850
rect 1498 1842 1514 1845
rect 1520 1851 1531 1853
rect 1520 1845 1522 1851
rect 1529 1845 1531 1851
rect 1520 1842 1531 1845
rect 372 1747 386 1749
rect 372 1740 374 1747
rect 382 1740 386 1747
rect 372 1734 386 1740
rect 393 1746 412 1749
rect 393 1737 396 1746
rect 406 1737 412 1746
rect 393 1734 412 1737
rect 431 1748 450 1749
rect 431 1740 437 1748
rect 445 1740 450 1748
rect 431 1734 450 1740
rect 457 1747 471 1749
rect 597 1754 614 1758
rect 457 1739 460 1747
rect 468 1739 471 1747
rect 457 1734 471 1739
rect 494 1747 513 1748
rect 494 1739 500 1747
rect 508 1739 513 1747
rect 494 1733 513 1739
rect 520 1746 534 1748
rect 520 1738 523 1746
rect 531 1738 534 1746
rect 597 1744 599 1754
rect 609 1744 614 1754
rect 597 1742 614 1744
rect 622 1755 637 1758
rect 622 1745 624 1755
rect 634 1745 637 1755
rect 622 1742 637 1745
rect 520 1733 534 1738
rect 295 1694 297 1703
rect 303 1694 305 1703
rect 313 1694 318 1703
rect 352 1588 366 1590
rect 352 1581 354 1588
rect 362 1581 366 1588
rect 352 1575 366 1581
rect 373 1587 392 1590
rect 373 1578 376 1587
rect 386 1578 392 1587
rect 373 1575 392 1578
rect 411 1589 430 1590
rect 411 1581 417 1589
rect 425 1581 430 1589
rect 411 1575 430 1581
rect 437 1588 451 1590
rect 437 1580 440 1588
rect 448 1580 451 1588
rect 437 1575 451 1580
rect 474 1588 493 1589
rect 474 1580 480 1588
rect 488 1580 493 1588
rect 474 1574 493 1580
rect 500 1587 514 1589
rect 617 1593 634 1597
rect 500 1579 503 1587
rect 511 1579 514 1587
rect 500 1574 514 1579
rect 542 1586 561 1587
rect 542 1578 548 1586
rect 556 1578 561 1586
rect 542 1572 561 1578
rect 568 1585 582 1587
rect 568 1577 571 1585
rect 579 1577 582 1585
rect 617 1583 619 1593
rect 629 1583 634 1593
rect 617 1581 634 1583
rect 642 1594 657 1597
rect 642 1584 644 1594
rect 654 1584 657 1594
rect 642 1581 657 1584
rect 568 1572 582 1577
rect 294 1539 296 1548
rect 302 1539 304 1548
rect 312 1539 317 1548
rect 361 1369 375 1371
rect 361 1362 363 1369
rect 371 1362 375 1369
rect 361 1356 375 1362
rect 382 1368 401 1371
rect 382 1359 385 1368
rect 395 1359 401 1368
rect 382 1356 401 1359
rect 420 1370 439 1371
rect 420 1362 426 1370
rect 434 1362 439 1370
rect 420 1356 439 1362
rect 446 1369 460 1371
rect 446 1361 449 1369
rect 457 1361 460 1369
rect 446 1356 460 1361
rect 483 1369 502 1370
rect 483 1361 489 1369
rect 497 1361 502 1369
rect 483 1355 502 1361
rect 509 1368 523 1370
rect 509 1360 512 1368
rect 520 1360 523 1368
rect 509 1355 523 1360
rect 551 1367 570 1368
rect 551 1359 557 1367
rect 565 1359 570 1367
rect 551 1353 570 1359
rect 577 1366 591 1368
rect 687 1373 704 1377
rect 577 1358 580 1366
rect 588 1358 591 1366
rect 577 1353 591 1358
rect 610 1366 629 1367
rect 610 1358 616 1366
rect 624 1358 629 1366
rect 610 1352 629 1358
rect 636 1365 650 1367
rect 636 1357 639 1365
rect 647 1357 650 1365
rect 687 1363 689 1373
rect 699 1363 704 1373
rect 687 1361 704 1363
rect 712 1374 727 1377
rect 712 1364 714 1374
rect 724 1364 727 1374
rect 712 1361 727 1364
rect 636 1352 650 1357
rect 294 1307 296 1316
rect 302 1307 304 1316
rect 312 1307 317 1316
rect 979 989 981 998
rect 987 989 989 998
rect 997 989 1002 998
rect 241 979 255 981
rect 241 972 243 979
rect 251 972 255 979
rect 241 966 255 972
rect 262 978 281 981
rect 262 969 265 978
rect 275 969 281 978
rect 262 966 281 969
rect 300 980 319 981
rect 300 972 306 980
rect 314 972 319 980
rect 300 966 319 972
rect 326 979 340 981
rect 326 971 329 979
rect 337 971 340 979
rect 326 966 340 971
rect 444 979 458 981
rect 444 972 446 979
rect 454 972 458 979
rect 444 966 458 972
rect 465 978 484 981
rect 465 969 468 978
rect 478 969 484 978
rect 465 966 484 969
rect 503 980 522 981
rect 503 972 509 980
rect 517 972 522 980
rect 503 966 522 972
rect 529 979 543 981
rect 529 971 532 979
rect 540 971 543 979
rect 529 966 543 971
rect 631 979 645 981
rect 631 972 633 979
rect 641 972 645 979
rect 631 966 645 972
rect 652 978 671 981
rect 652 969 655 978
rect 665 969 671 978
rect 652 966 671 969
rect 690 980 709 981
rect 690 972 696 980
rect 704 972 709 980
rect 690 966 709 972
rect 716 979 730 981
rect 716 971 719 979
rect 727 971 730 979
rect 716 966 730 971
rect 812 979 826 981
rect 812 972 814 979
rect 822 972 826 979
rect 812 966 826 972
rect 833 978 852 981
rect 833 969 836 978
rect 846 969 852 978
rect 833 966 852 969
rect 871 980 890 981
rect 871 972 877 980
rect 885 972 890 980
rect 871 966 890 972
rect 897 979 911 981
rect 897 971 900 979
rect 908 971 911 979
rect 897 966 911 971
rect 981 697 983 706
rect 989 697 991 706
rect 999 697 1004 706
rect 247 690 261 692
rect 247 683 249 690
rect 257 683 261 690
rect 247 677 261 683
rect 268 689 287 692
rect 268 680 271 689
rect 281 680 287 689
rect 268 677 287 680
rect 306 691 325 692
rect 306 683 312 691
rect 320 683 325 691
rect 306 677 325 683
rect 332 690 346 692
rect 332 682 335 690
rect 343 682 346 690
rect 332 677 346 682
rect 450 690 464 692
rect 450 683 452 690
rect 460 683 464 690
rect 450 677 464 683
rect 471 689 490 692
rect 471 680 474 689
rect 484 680 490 689
rect 471 677 490 680
rect 509 691 528 692
rect 509 683 515 691
rect 523 683 528 691
rect 509 677 528 683
rect 535 690 549 692
rect 535 682 538 690
rect 546 682 549 690
rect 535 677 549 682
rect 637 690 651 692
rect 637 683 639 690
rect 647 683 651 690
rect 637 677 651 683
rect 658 689 677 692
rect 658 680 661 689
rect 671 680 677 689
rect 658 677 677 680
rect 696 691 715 692
rect 696 683 702 691
rect 710 683 715 691
rect 696 677 715 683
rect 722 690 736 692
rect 722 682 725 690
rect 733 682 736 690
rect 722 677 736 682
rect 818 690 832 692
rect 818 683 820 690
rect 828 683 832 690
rect 818 677 832 683
rect 839 689 858 692
rect 839 680 842 689
rect 852 680 858 689
rect 839 677 858 680
rect 877 691 896 692
rect 877 683 883 691
rect 891 683 896 691
rect 877 677 896 683
rect 903 690 917 692
rect 903 682 906 690
rect 914 682 917 690
rect 903 677 917 682
rect 1006 380 1008 389
rect 1014 380 1016 389
rect 1024 380 1029 389
rect 267 373 281 375
rect 267 366 269 373
rect 277 366 281 373
rect 267 360 281 366
rect 288 372 307 375
rect 288 363 291 372
rect 301 363 307 372
rect 288 360 307 363
rect 326 374 345 375
rect 326 366 332 374
rect 340 366 345 374
rect 326 360 345 366
rect 352 373 366 375
rect 352 365 355 373
rect 363 365 366 373
rect 352 360 366 365
rect 470 373 484 375
rect 470 366 472 373
rect 480 366 484 373
rect 470 360 484 366
rect 491 372 510 375
rect 491 363 494 372
rect 504 363 510 372
rect 491 360 510 363
rect 529 374 548 375
rect 529 366 535 374
rect 543 366 548 374
rect 529 360 548 366
rect 555 373 569 375
rect 555 365 558 373
rect 566 365 569 373
rect 555 360 569 365
rect 657 373 671 375
rect 657 366 659 373
rect 667 366 671 373
rect 657 360 671 366
rect 678 372 697 375
rect 678 363 681 372
rect 691 363 697 372
rect 678 360 697 363
rect 716 374 735 375
rect 716 366 722 374
rect 730 366 735 374
rect 716 360 735 366
rect 742 373 756 375
rect 742 365 745 373
rect 753 365 756 373
rect 742 360 756 365
rect 838 373 852 375
rect 838 366 840 373
rect 848 366 852 373
rect 838 360 852 366
rect 859 372 878 375
rect 859 363 862 372
rect 872 363 878 372
rect 859 360 878 363
rect 897 374 916 375
rect 897 366 903 374
rect 911 366 916 374
rect 897 360 916 366
rect 923 373 937 375
rect 923 365 926 373
rect 934 365 937 373
rect 923 360 937 365
rect 1015 89 1017 98
rect 1023 89 1025 98
rect 1033 89 1038 98
rect 265 82 279 84
rect 265 75 267 82
rect 275 75 279 82
rect 265 69 279 75
rect 286 81 305 84
rect 286 72 289 81
rect 299 72 305 81
rect 286 69 305 72
rect 324 83 343 84
rect 324 75 330 83
rect 338 75 343 83
rect 324 69 343 75
rect 350 82 364 84
rect 350 74 353 82
rect 361 74 364 82
rect 350 69 364 74
rect 468 82 482 84
rect 468 75 470 82
rect 478 75 482 82
rect 468 69 482 75
rect 489 81 508 84
rect 489 72 492 81
rect 502 72 508 81
rect 489 69 508 72
rect 527 83 546 84
rect 527 75 533 83
rect 541 75 546 83
rect 527 69 546 75
rect 553 82 567 84
rect 553 74 556 82
rect 564 74 567 82
rect 553 69 567 74
rect 655 82 669 84
rect 655 75 657 82
rect 665 75 669 82
rect 655 69 669 75
rect 676 81 695 84
rect 676 72 679 81
rect 689 72 695 81
rect 676 69 695 72
rect 714 83 733 84
rect 714 75 720 83
rect 728 75 733 83
rect 714 69 733 75
rect 740 82 754 84
rect 740 74 743 82
rect 751 74 754 82
rect 740 69 754 74
rect 836 82 850 84
rect 836 75 838 82
rect 846 75 850 82
rect 836 69 850 75
rect 857 81 876 84
rect 857 72 860 81
rect 870 72 876 81
rect 857 69 876 72
rect 895 83 914 84
rect 895 75 901 83
rect 909 75 914 83
rect 895 69 914 75
rect 921 82 935 84
rect 921 74 924 82
rect 932 74 935 82
rect 921 69 935 74
rect 318 -350 332 -348
rect 318 -357 320 -350
rect 328 -357 332 -350
rect 318 -363 332 -357
rect 339 -351 358 -348
rect 339 -360 342 -351
rect 352 -360 358 -351
rect 339 -363 358 -360
rect 377 -349 396 -348
rect 377 -357 383 -349
rect 391 -357 396 -349
rect 377 -363 396 -357
rect 403 -350 417 -348
rect 403 -358 406 -350
rect 414 -358 417 -350
rect 403 -363 417 -358
rect 488 -357 505 -353
rect 488 -367 490 -357
rect 500 -367 505 -357
rect 488 -369 505 -367
rect 513 -356 528 -353
rect 513 -366 515 -356
rect 525 -366 528 -356
rect 513 -369 528 -366
rect 239 -410 241 -401
rect 247 -410 249 -401
rect 257 -410 262 -401
rect 318 -519 332 -517
rect 318 -526 320 -519
rect 328 -526 332 -519
rect 318 -532 332 -526
rect 339 -520 358 -517
rect 339 -529 342 -520
rect 352 -529 358 -520
rect 339 -532 358 -529
rect 377 -518 396 -517
rect 377 -526 383 -518
rect 391 -526 396 -518
rect 377 -532 396 -526
rect 403 -519 417 -517
rect 543 -512 560 -508
rect 403 -527 406 -519
rect 414 -527 417 -519
rect 403 -532 417 -527
rect 440 -519 459 -518
rect 440 -527 446 -519
rect 454 -527 459 -519
rect 440 -533 459 -527
rect 466 -520 480 -518
rect 466 -528 469 -520
rect 477 -528 480 -520
rect 543 -522 545 -512
rect 555 -522 560 -512
rect 543 -524 560 -522
rect 568 -511 583 -508
rect 568 -521 570 -511
rect 580 -521 583 -511
rect 568 -524 583 -521
rect 466 -533 480 -528
rect 1468 416 1470 425
rect 1476 416 1478 425
rect 1486 416 1491 425
rect 1190 405 1204 407
rect 1190 398 1192 405
rect 1200 398 1204 405
rect 1190 392 1204 398
rect 1211 404 1230 407
rect 1211 395 1214 404
rect 1224 395 1230 404
rect 1211 392 1230 395
rect 1249 406 1268 407
rect 1249 398 1255 406
rect 1263 398 1268 406
rect 1249 392 1268 398
rect 1275 405 1289 407
rect 1275 397 1278 405
rect 1286 397 1289 405
rect 1275 392 1289 397
rect 1325 406 1341 408
rect 1325 398 1331 406
rect 1339 398 1341 406
rect 1325 393 1341 398
rect 1348 405 1367 408
rect 1348 396 1351 405
rect 1361 396 1367 405
rect 1348 393 1367 396
rect 1386 407 1405 408
rect 1386 399 1392 407
rect 1400 399 1405 407
rect 1386 393 1405 399
rect 1412 406 1426 408
rect 1412 398 1415 406
rect 1423 398 1426 406
rect 1412 393 1426 398
rect 241 -572 243 -563
rect 249 -572 251 -563
rect 259 -572 264 -563
rect 298 -678 312 -676
rect 298 -685 300 -678
rect 308 -685 312 -678
rect 298 -691 312 -685
rect 319 -679 338 -676
rect 319 -688 322 -679
rect 332 -688 338 -679
rect 319 -691 338 -688
rect 357 -677 376 -676
rect 357 -685 363 -677
rect 371 -685 376 -677
rect 357 -691 376 -685
rect 383 -678 397 -676
rect 383 -686 386 -678
rect 394 -686 397 -678
rect 383 -691 397 -686
rect 420 -678 439 -677
rect 420 -686 426 -678
rect 434 -686 439 -678
rect 420 -692 439 -686
rect 446 -679 460 -677
rect 563 -673 580 -669
rect 446 -687 449 -679
rect 457 -687 460 -679
rect 446 -692 460 -687
rect 488 -680 507 -679
rect 488 -688 494 -680
rect 502 -688 507 -680
rect 488 -694 507 -688
rect 514 -681 528 -679
rect 514 -689 517 -681
rect 525 -689 528 -681
rect 563 -683 565 -673
rect 575 -683 580 -673
rect 563 -685 580 -683
rect 588 -672 603 -669
rect 588 -682 590 -672
rect 600 -682 603 -672
rect 588 -685 603 -682
rect 514 -694 528 -689
rect 240 -727 242 -718
rect 248 -727 250 -718
rect 258 -727 263 -718
rect 307 -897 321 -895
rect 307 -904 309 -897
rect 317 -904 321 -897
rect 307 -910 321 -904
rect 328 -898 347 -895
rect 328 -907 331 -898
rect 341 -907 347 -898
rect 328 -910 347 -907
rect 366 -896 385 -895
rect 366 -904 372 -896
rect 380 -904 385 -896
rect 366 -910 385 -904
rect 392 -897 406 -895
rect 392 -905 395 -897
rect 403 -905 406 -897
rect 392 -910 406 -905
rect 429 -897 448 -896
rect 429 -905 435 -897
rect 443 -905 448 -897
rect 429 -911 448 -905
rect 455 -898 469 -896
rect 455 -906 458 -898
rect 466 -906 469 -898
rect 455 -911 469 -906
rect 497 -899 516 -898
rect 497 -907 503 -899
rect 511 -907 516 -899
rect 497 -913 516 -907
rect 523 -900 537 -898
rect 633 -893 650 -889
rect 523 -908 526 -900
rect 534 -908 537 -900
rect 523 -913 537 -908
rect 556 -900 575 -899
rect 556 -908 562 -900
rect 570 -908 575 -900
rect 556 -914 575 -908
rect 582 -901 596 -899
rect 582 -909 585 -901
rect 593 -909 596 -901
rect 633 -903 635 -893
rect 645 -903 650 -893
rect 633 -905 650 -903
rect 658 -892 673 -889
rect 658 -902 660 -892
rect 670 -902 673 -892
rect 658 -905 673 -902
rect 582 -914 596 -909
rect 1398 -416 1409 -413
rect 1398 -421 1400 -416
rect 1406 -421 1409 -416
rect 1398 -424 1409 -421
rect 1415 -415 1431 -413
rect 1415 -421 1419 -415
rect 1426 -421 1431 -415
rect 1415 -424 1431 -421
rect 1436 -416 1450 -413
rect 1436 -421 1440 -416
rect 1446 -421 1450 -416
rect 1436 -424 1450 -421
rect 1456 -415 1469 -413
rect 1456 -421 1459 -415
rect 1466 -421 1469 -415
rect 1456 -424 1469 -421
rect 1475 -416 1489 -413
rect 1475 -422 1479 -416
rect 1485 -422 1489 -416
rect 1475 -424 1489 -422
rect 1495 -414 1508 -413
rect 1495 -421 1498 -414
rect 1505 -421 1508 -414
rect 1495 -424 1508 -421
rect 1518 -416 1532 -413
rect 1518 -422 1522 -416
rect 1528 -422 1532 -416
rect 1518 -424 1532 -422
rect 1538 -415 1551 -413
rect 1538 -421 1540 -415
rect 1547 -421 1551 -415
rect 1538 -424 1551 -421
rect 1558 -416 1574 -413
rect 1558 -421 1564 -416
rect 1570 -421 1574 -416
rect 1558 -424 1574 -421
rect 1580 -415 1591 -413
rect 1580 -421 1582 -415
rect 1589 -421 1591 -415
rect 1580 -424 1591 -421
rect 240 -959 242 -950
rect 248 -959 250 -950
rect 258 -959 263 -950
<< pdiffusion >>
rect 372 2001 386 2003
rect 372 1995 375 2001
rect 382 1995 386 2001
rect 372 1988 386 1995
rect 393 1999 412 2003
rect 393 1991 397 1999
rect 406 1991 412 1999
rect 393 1988 412 1991
rect 439 1999 450 2003
rect 439 1992 441 1999
rect 449 1992 450 1999
rect 439 1988 450 1992
rect 457 1997 479 2003
rect 457 1991 460 1997
rect 468 1991 479 1997
rect 457 1988 479 1991
rect 543 1981 545 1991
rect 555 1981 559 1991
rect 543 1975 559 1981
rect 567 1988 583 1991
rect 567 1978 569 1988
rect 579 1978 583 1988
rect 567 1975 583 1978
rect 293 1907 295 1916
rect 301 1907 303 1916
rect 312 1907 316 1916
rect 1338 1912 1349 1914
rect 1338 1906 1340 1912
rect 1346 1906 1349 1912
rect 1338 1903 1349 1906
rect 1355 1909 1371 1914
rect 1355 1903 1359 1909
rect 1365 1903 1371 1909
rect 1376 1909 1390 1914
rect 1376 1903 1380 1909
rect 1386 1903 1390 1909
rect 1396 1909 1409 1914
rect 1396 1903 1400 1909
rect 1406 1903 1409 1909
rect 1415 1909 1429 1914
rect 1415 1903 1419 1909
rect 1425 1903 1429 1909
rect 1435 1909 1448 1914
rect 1435 1903 1438 1909
rect 1444 1903 1448 1909
rect 1458 1909 1472 1914
rect 1458 1903 1462 1909
rect 1468 1903 1472 1909
rect 1478 1909 1491 1914
rect 1478 1903 1481 1909
rect 1487 1903 1491 1909
rect 1501 1912 1514 1914
rect 1501 1906 1504 1912
rect 1510 1906 1514 1912
rect 1501 1903 1514 1906
rect 1520 1910 1534 1914
rect 1520 1904 1522 1910
rect 1529 1904 1534 1910
rect 1520 1903 1534 1904
rect 372 1832 386 1834
rect 372 1826 375 1832
rect 382 1826 386 1832
rect 372 1819 386 1826
rect 393 1830 412 1834
rect 393 1822 397 1830
rect 406 1822 412 1830
rect 393 1819 412 1822
rect 439 1830 450 1834
rect 439 1823 441 1830
rect 449 1823 450 1830
rect 439 1819 450 1823
rect 457 1828 479 1834
rect 457 1822 460 1828
rect 468 1822 479 1828
rect 457 1819 479 1822
rect 502 1829 513 1833
rect 502 1822 504 1829
rect 512 1822 513 1829
rect 295 1745 297 1754
rect 303 1745 305 1754
rect 314 1745 318 1754
rect 502 1818 513 1822
rect 520 1827 542 1833
rect 520 1821 523 1827
rect 531 1821 542 1827
rect 520 1818 542 1821
rect 598 1826 600 1836
rect 610 1826 614 1836
rect 598 1820 614 1826
rect 622 1833 638 1836
rect 622 1823 624 1833
rect 634 1823 638 1833
rect 622 1820 638 1823
rect 352 1673 366 1675
rect 352 1667 355 1673
rect 362 1667 366 1673
rect 352 1660 366 1667
rect 373 1671 392 1675
rect 373 1663 377 1671
rect 386 1663 392 1671
rect 373 1660 392 1663
rect 419 1671 430 1675
rect 419 1664 421 1671
rect 429 1664 430 1671
rect 419 1660 430 1664
rect 437 1669 459 1675
rect 437 1663 440 1669
rect 448 1663 459 1669
rect 437 1660 459 1663
rect 482 1670 493 1674
rect 482 1663 484 1670
rect 492 1663 493 1670
rect 294 1590 296 1599
rect 302 1590 304 1599
rect 313 1590 317 1599
rect 482 1659 493 1663
rect 500 1668 522 1674
rect 500 1662 503 1668
rect 511 1662 522 1668
rect 500 1659 522 1662
rect 550 1668 561 1672
rect 550 1661 552 1668
rect 560 1661 561 1668
rect 550 1657 561 1661
rect 568 1666 590 1672
rect 568 1660 571 1666
rect 579 1660 590 1666
rect 568 1657 590 1660
rect 618 1665 620 1675
rect 630 1665 634 1675
rect 618 1659 634 1665
rect 642 1672 658 1675
rect 642 1662 644 1672
rect 654 1662 658 1672
rect 642 1659 658 1662
rect 361 1454 375 1456
rect 361 1448 364 1454
rect 371 1448 375 1454
rect 361 1441 375 1448
rect 382 1452 401 1456
rect 382 1444 386 1452
rect 395 1444 401 1452
rect 382 1441 401 1444
rect 428 1452 439 1456
rect 428 1445 430 1452
rect 438 1445 439 1452
rect 428 1441 439 1445
rect 446 1450 468 1456
rect 446 1444 449 1450
rect 457 1444 468 1450
rect 446 1441 468 1444
rect 491 1451 502 1455
rect 491 1444 493 1451
rect 501 1444 502 1451
rect 491 1440 502 1444
rect 509 1449 531 1455
rect 509 1443 512 1449
rect 520 1443 531 1449
rect 509 1440 531 1443
rect 559 1449 570 1453
rect 559 1442 561 1449
rect 569 1442 570 1449
rect 294 1358 296 1367
rect 302 1358 304 1367
rect 313 1358 317 1367
rect 559 1438 570 1442
rect 577 1447 599 1453
rect 577 1441 580 1447
rect 588 1441 599 1447
rect 577 1438 599 1441
rect 618 1448 629 1452
rect 618 1441 620 1448
rect 628 1441 629 1448
rect 618 1437 629 1441
rect 636 1446 658 1452
rect 636 1440 639 1446
rect 647 1440 658 1446
rect 636 1437 658 1440
rect 688 1445 690 1455
rect 700 1445 704 1455
rect 688 1439 704 1445
rect 712 1452 728 1455
rect 712 1442 714 1452
rect 724 1442 728 1452
rect 712 1439 728 1442
rect 241 1064 255 1066
rect 241 1058 244 1064
rect 251 1058 255 1064
rect 241 1051 255 1058
rect 262 1062 281 1066
rect 262 1054 266 1062
rect 275 1054 281 1062
rect 262 1051 281 1054
rect 308 1062 319 1066
rect 308 1055 310 1062
rect 318 1055 319 1062
rect 308 1051 319 1055
rect 326 1060 348 1066
rect 326 1054 329 1060
rect 337 1054 348 1060
rect 326 1051 348 1054
rect 444 1064 458 1066
rect 444 1058 447 1064
rect 454 1058 458 1064
rect 444 1051 458 1058
rect 465 1062 484 1066
rect 465 1054 469 1062
rect 478 1054 484 1062
rect 465 1051 484 1054
rect 511 1062 522 1066
rect 511 1055 513 1062
rect 521 1055 522 1062
rect 511 1051 522 1055
rect 529 1060 551 1066
rect 529 1054 532 1060
rect 540 1054 551 1060
rect 529 1051 551 1054
rect 631 1064 645 1066
rect 631 1058 634 1064
rect 641 1058 645 1064
rect 631 1051 645 1058
rect 652 1062 671 1066
rect 652 1054 656 1062
rect 665 1054 671 1062
rect 652 1051 671 1054
rect 698 1062 709 1066
rect 698 1055 700 1062
rect 708 1055 709 1062
rect 698 1051 709 1055
rect 716 1060 738 1066
rect 716 1054 719 1060
rect 727 1054 738 1060
rect 716 1051 738 1054
rect 812 1064 826 1066
rect 812 1058 815 1064
rect 822 1058 826 1064
rect 812 1051 826 1058
rect 833 1062 852 1066
rect 833 1054 837 1062
rect 846 1054 852 1062
rect 833 1051 852 1054
rect 879 1062 890 1066
rect 879 1055 881 1062
rect 889 1055 890 1062
rect 879 1051 890 1055
rect 897 1060 919 1066
rect 897 1054 900 1060
rect 908 1054 919 1060
rect 897 1051 919 1054
rect 979 1040 981 1049
rect 987 1040 989 1049
rect 998 1040 1002 1049
rect 247 775 261 777
rect 247 769 250 775
rect 257 769 261 775
rect 247 762 261 769
rect 268 773 287 777
rect 268 765 272 773
rect 281 765 287 773
rect 268 762 287 765
rect 314 773 325 777
rect 314 766 316 773
rect 324 766 325 773
rect 314 762 325 766
rect 332 771 354 777
rect 332 765 335 771
rect 343 765 354 771
rect 332 762 354 765
rect 450 775 464 777
rect 450 769 453 775
rect 460 769 464 775
rect 450 762 464 769
rect 471 773 490 777
rect 471 765 475 773
rect 484 765 490 773
rect 471 762 490 765
rect 517 773 528 777
rect 517 766 519 773
rect 527 766 528 773
rect 517 762 528 766
rect 535 771 557 777
rect 535 765 538 771
rect 546 765 557 771
rect 535 762 557 765
rect 637 775 651 777
rect 637 769 640 775
rect 647 769 651 775
rect 637 762 651 769
rect 658 773 677 777
rect 658 765 662 773
rect 671 765 677 773
rect 658 762 677 765
rect 704 773 715 777
rect 704 766 706 773
rect 714 766 715 773
rect 704 762 715 766
rect 722 771 744 777
rect 722 765 725 771
rect 733 765 744 771
rect 722 762 744 765
rect 818 775 832 777
rect 818 769 821 775
rect 828 769 832 775
rect 818 762 832 769
rect 839 773 858 777
rect 839 765 843 773
rect 852 765 858 773
rect 839 762 858 765
rect 885 773 896 777
rect 885 766 887 773
rect 895 766 896 773
rect 885 762 896 766
rect 903 771 925 777
rect 903 765 906 771
rect 914 765 925 771
rect 903 762 925 765
rect 981 748 983 757
rect 989 748 991 757
rect 1000 748 1004 757
rect 267 458 281 460
rect 267 452 270 458
rect 277 452 281 458
rect 267 445 281 452
rect 288 456 307 460
rect 288 448 292 456
rect 301 448 307 456
rect 288 445 307 448
rect 334 456 345 460
rect 334 449 336 456
rect 344 449 345 456
rect 334 445 345 449
rect 352 454 374 460
rect 352 448 355 454
rect 363 448 374 454
rect 352 445 374 448
rect 470 458 484 460
rect 470 452 473 458
rect 480 452 484 458
rect 470 445 484 452
rect 491 456 510 460
rect 491 448 495 456
rect 504 448 510 456
rect 491 445 510 448
rect 537 456 548 460
rect 537 449 539 456
rect 547 449 548 456
rect 537 445 548 449
rect 555 454 577 460
rect 555 448 558 454
rect 566 448 577 454
rect 555 445 577 448
rect 657 458 671 460
rect 657 452 660 458
rect 667 452 671 458
rect 657 445 671 452
rect 678 456 697 460
rect 678 448 682 456
rect 691 448 697 456
rect 678 445 697 448
rect 724 456 735 460
rect 724 449 726 456
rect 734 449 735 456
rect 724 445 735 449
rect 742 454 764 460
rect 742 448 745 454
rect 753 448 764 454
rect 742 445 764 448
rect 838 458 852 460
rect 838 452 841 458
rect 848 452 852 458
rect 838 445 852 452
rect 859 456 878 460
rect 859 448 863 456
rect 872 448 878 456
rect 859 445 878 448
rect 905 456 916 460
rect 905 449 907 456
rect 915 449 916 456
rect 905 445 916 449
rect 923 454 945 460
rect 923 448 926 454
rect 934 448 945 454
rect 923 445 945 448
rect 1006 431 1008 440
rect 1014 431 1016 440
rect 1025 431 1029 440
rect 265 167 279 169
rect 265 161 268 167
rect 275 161 279 167
rect 265 154 279 161
rect 286 165 305 169
rect 286 157 290 165
rect 299 157 305 165
rect 286 154 305 157
rect 332 165 343 169
rect 332 158 334 165
rect 342 158 343 165
rect 332 154 343 158
rect 350 163 372 169
rect 350 157 353 163
rect 361 157 372 163
rect 350 154 372 157
rect 468 167 482 169
rect 468 161 471 167
rect 478 161 482 167
rect 468 154 482 161
rect 489 165 508 169
rect 489 157 493 165
rect 502 157 508 165
rect 489 154 508 157
rect 535 165 546 169
rect 535 158 537 165
rect 545 158 546 165
rect 535 154 546 158
rect 553 163 575 169
rect 553 157 556 163
rect 564 157 575 163
rect 553 154 575 157
rect 655 167 669 169
rect 655 161 658 167
rect 665 161 669 167
rect 655 154 669 161
rect 676 165 695 169
rect 676 157 680 165
rect 689 157 695 165
rect 676 154 695 157
rect 722 165 733 169
rect 722 158 724 165
rect 732 158 733 165
rect 722 154 733 158
rect 740 163 762 169
rect 740 157 743 163
rect 751 157 762 163
rect 740 154 762 157
rect 836 167 850 169
rect 836 161 839 167
rect 846 161 850 167
rect 836 154 850 161
rect 857 165 876 169
rect 857 157 861 165
rect 870 157 876 165
rect 857 154 876 157
rect 903 165 914 169
rect 903 158 905 165
rect 913 158 914 165
rect 903 154 914 158
rect 921 163 943 169
rect 921 157 924 163
rect 932 157 943 163
rect 921 154 943 157
rect 1015 140 1017 149
rect 1023 140 1025 149
rect 1034 140 1038 149
rect 318 -265 332 -263
rect 318 -271 321 -265
rect 328 -271 332 -265
rect 318 -278 332 -271
rect 339 -267 358 -263
rect 339 -275 343 -267
rect 352 -275 358 -267
rect 339 -278 358 -275
rect 385 -267 396 -263
rect 385 -274 387 -267
rect 395 -274 396 -267
rect 385 -278 396 -274
rect 403 -269 425 -263
rect 403 -275 406 -269
rect 414 -275 425 -269
rect 403 -278 425 -275
rect 489 -285 491 -275
rect 501 -285 505 -275
rect 489 -291 505 -285
rect 513 -278 529 -275
rect 513 -288 515 -278
rect 525 -288 529 -278
rect 513 -291 529 -288
rect 239 -359 241 -350
rect 247 -359 249 -350
rect 258 -359 262 -350
rect 318 -434 332 -432
rect 318 -440 321 -434
rect 328 -440 332 -434
rect 318 -447 332 -440
rect 339 -436 358 -432
rect 339 -444 343 -436
rect 352 -444 358 -436
rect 339 -447 358 -444
rect 385 -436 396 -432
rect 385 -443 387 -436
rect 395 -443 396 -436
rect 385 -447 396 -443
rect 403 -438 425 -432
rect 403 -444 406 -438
rect 414 -444 425 -438
rect 403 -447 425 -444
rect 448 -437 459 -433
rect 448 -444 450 -437
rect 458 -444 459 -437
rect 241 -521 243 -512
rect 249 -521 251 -512
rect 260 -521 264 -512
rect 448 -448 459 -444
rect 466 -439 488 -433
rect 466 -445 469 -439
rect 477 -445 488 -439
rect 466 -448 488 -445
rect 544 -440 546 -430
rect 556 -440 560 -430
rect 544 -446 560 -440
rect 568 -433 584 -430
rect 568 -443 570 -433
rect 580 -443 584 -433
rect 568 -446 584 -443
rect 1190 490 1204 492
rect 1190 484 1193 490
rect 1200 484 1204 490
rect 1190 477 1204 484
rect 1211 488 1230 492
rect 1211 480 1215 488
rect 1224 480 1230 488
rect 1211 477 1230 480
rect 1257 488 1268 492
rect 1257 481 1259 488
rect 1267 481 1268 488
rect 1257 477 1268 481
rect 1275 486 1297 492
rect 1275 480 1278 486
rect 1286 480 1297 486
rect 1275 477 1297 480
rect 1327 491 1341 493
rect 1327 485 1330 491
rect 1337 485 1341 491
rect 1327 478 1341 485
rect 1348 489 1367 493
rect 1348 481 1352 489
rect 1361 481 1367 489
rect 1348 478 1367 481
rect 1394 489 1405 493
rect 1394 482 1396 489
rect 1404 482 1405 489
rect 1394 478 1405 482
rect 1412 487 1434 493
rect 1412 481 1415 487
rect 1423 481 1434 487
rect 1412 478 1434 481
rect 1468 467 1470 476
rect 1476 467 1478 476
rect 1487 467 1491 476
rect 298 -593 312 -591
rect 298 -599 301 -593
rect 308 -599 312 -593
rect 298 -606 312 -599
rect 319 -595 338 -591
rect 319 -603 323 -595
rect 332 -603 338 -595
rect 319 -606 338 -603
rect 365 -595 376 -591
rect 365 -602 367 -595
rect 375 -602 376 -595
rect 365 -606 376 -602
rect 383 -597 405 -591
rect 383 -603 386 -597
rect 394 -603 405 -597
rect 383 -606 405 -603
rect 428 -596 439 -592
rect 428 -603 430 -596
rect 438 -603 439 -596
rect 240 -676 242 -667
rect 248 -676 250 -667
rect 259 -676 263 -667
rect 428 -607 439 -603
rect 446 -598 468 -592
rect 446 -604 449 -598
rect 457 -604 468 -598
rect 446 -607 468 -604
rect 496 -598 507 -594
rect 496 -605 498 -598
rect 506 -605 507 -598
rect 496 -609 507 -605
rect 514 -600 536 -594
rect 514 -606 517 -600
rect 525 -606 536 -600
rect 514 -609 536 -606
rect 564 -601 566 -591
rect 576 -601 580 -591
rect 564 -607 580 -601
rect 588 -594 604 -591
rect 588 -604 590 -594
rect 600 -604 604 -594
rect 588 -607 604 -604
rect 307 -812 321 -810
rect 307 -818 310 -812
rect 317 -818 321 -812
rect 307 -825 321 -818
rect 328 -814 347 -810
rect 328 -822 332 -814
rect 341 -822 347 -814
rect 328 -825 347 -822
rect 374 -814 385 -810
rect 374 -821 376 -814
rect 384 -821 385 -814
rect 374 -825 385 -821
rect 392 -816 414 -810
rect 392 -822 395 -816
rect 403 -822 414 -816
rect 392 -825 414 -822
rect 437 -815 448 -811
rect 437 -822 439 -815
rect 447 -822 448 -815
rect 437 -826 448 -822
rect 455 -817 477 -811
rect 455 -823 458 -817
rect 466 -823 477 -817
rect 455 -826 477 -823
rect 505 -817 516 -813
rect 505 -824 507 -817
rect 515 -824 516 -817
rect 240 -908 242 -899
rect 248 -908 250 -899
rect 259 -908 263 -899
rect 505 -828 516 -824
rect 523 -819 545 -813
rect 523 -825 526 -819
rect 534 -825 545 -819
rect 523 -828 545 -825
rect 564 -818 575 -814
rect 564 -825 566 -818
rect 574 -825 575 -818
rect 564 -829 575 -825
rect 582 -820 604 -814
rect 582 -826 585 -820
rect 593 -826 604 -820
rect 582 -829 604 -826
rect 634 -821 636 -811
rect 646 -821 650 -811
rect 634 -827 650 -821
rect 658 -814 674 -811
rect 658 -824 660 -814
rect 670 -824 674 -814
rect 658 -827 674 -824
rect 1398 -354 1409 -352
rect 1398 -360 1400 -354
rect 1406 -360 1409 -354
rect 1398 -363 1409 -360
rect 1415 -357 1431 -352
rect 1415 -363 1419 -357
rect 1425 -363 1431 -357
rect 1436 -357 1450 -352
rect 1436 -363 1440 -357
rect 1446 -363 1450 -357
rect 1456 -357 1469 -352
rect 1456 -363 1460 -357
rect 1466 -363 1469 -357
rect 1475 -357 1489 -352
rect 1475 -363 1479 -357
rect 1485 -363 1489 -357
rect 1495 -357 1508 -352
rect 1495 -363 1498 -357
rect 1504 -363 1508 -357
rect 1518 -357 1532 -352
rect 1518 -363 1522 -357
rect 1528 -363 1532 -357
rect 1538 -357 1551 -352
rect 1538 -363 1541 -357
rect 1547 -363 1551 -357
rect 1561 -354 1574 -352
rect 1561 -360 1564 -354
rect 1570 -360 1574 -354
rect 1561 -363 1574 -360
rect 1580 -356 1594 -352
rect 1580 -362 1582 -356
rect 1589 -362 1594 -356
rect 1580 -363 1594 -362
<< ndcontact >>
rect 374 1909 382 1916
rect 396 1906 406 1915
rect 437 1909 445 1917
rect 460 1908 468 1916
rect 544 1899 554 1909
rect 569 1900 579 1910
rect 285 1856 293 1865
rect 303 1856 311 1865
rect 1340 1845 1346 1850
rect 1359 1845 1366 1851
rect 1380 1845 1386 1850
rect 1399 1845 1406 1851
rect 1419 1844 1425 1850
rect 1438 1845 1445 1852
rect 1462 1844 1468 1850
rect 1480 1845 1487 1851
rect 1504 1845 1510 1850
rect 1522 1845 1529 1851
rect 374 1740 382 1747
rect 396 1737 406 1746
rect 437 1740 445 1748
rect 460 1739 468 1747
rect 500 1739 508 1747
rect 523 1738 531 1746
rect 599 1744 609 1754
rect 624 1745 634 1755
rect 287 1694 295 1703
rect 305 1694 313 1703
rect 354 1581 362 1588
rect 376 1578 386 1587
rect 417 1581 425 1589
rect 440 1580 448 1588
rect 480 1580 488 1588
rect 503 1579 511 1587
rect 548 1578 556 1586
rect 571 1577 579 1585
rect 619 1583 629 1593
rect 644 1584 654 1594
rect 286 1539 294 1548
rect 304 1539 312 1548
rect 363 1362 371 1369
rect 385 1359 395 1368
rect 426 1362 434 1370
rect 449 1361 457 1369
rect 489 1361 497 1369
rect 512 1360 520 1368
rect 557 1359 565 1367
rect 580 1358 588 1366
rect 616 1358 624 1366
rect 639 1357 647 1365
rect 689 1363 699 1373
rect 714 1364 724 1374
rect 286 1307 294 1316
rect 304 1307 312 1316
rect 971 989 979 998
rect 989 989 997 998
rect 243 972 251 979
rect 265 969 275 978
rect 306 972 314 980
rect 329 971 337 979
rect 446 972 454 979
rect 468 969 478 978
rect 509 972 517 980
rect 532 971 540 979
rect 633 972 641 979
rect 655 969 665 978
rect 696 972 704 980
rect 719 971 727 979
rect 814 972 822 979
rect 836 969 846 978
rect 877 972 885 980
rect 900 971 908 979
rect 973 697 981 706
rect 991 697 999 706
rect 249 683 257 690
rect 271 680 281 689
rect 312 683 320 691
rect 335 682 343 690
rect 452 683 460 690
rect 474 680 484 689
rect 515 683 523 691
rect 538 682 546 690
rect 639 683 647 690
rect 661 680 671 689
rect 702 683 710 691
rect 725 682 733 690
rect 820 683 828 690
rect 842 680 852 689
rect 883 683 891 691
rect 906 682 914 690
rect 998 380 1006 389
rect 1016 380 1024 389
rect 269 366 277 373
rect 291 363 301 372
rect 332 366 340 374
rect 355 365 363 373
rect 472 366 480 373
rect 494 363 504 372
rect 535 366 543 374
rect 558 365 566 373
rect 659 366 667 373
rect 681 363 691 372
rect 722 366 730 374
rect 745 365 753 373
rect 840 366 848 373
rect 862 363 872 372
rect 903 366 911 374
rect 926 365 934 373
rect 1007 89 1015 98
rect 1025 89 1033 98
rect 267 75 275 82
rect 289 72 299 81
rect 330 75 338 83
rect 353 74 361 82
rect 470 75 478 82
rect 492 72 502 81
rect 533 75 541 83
rect 556 74 564 82
rect 657 75 665 82
rect 679 72 689 81
rect 720 75 728 83
rect 743 74 751 82
rect 838 75 846 82
rect 860 72 870 81
rect 901 75 909 83
rect 924 74 932 82
rect 320 -357 328 -350
rect 342 -360 352 -351
rect 383 -357 391 -349
rect 406 -358 414 -350
rect 490 -367 500 -357
rect 515 -366 525 -356
rect 231 -410 239 -401
rect 249 -410 257 -401
rect 320 -526 328 -519
rect 342 -529 352 -520
rect 383 -526 391 -518
rect 406 -527 414 -519
rect 446 -527 454 -519
rect 469 -528 477 -520
rect 545 -522 555 -512
rect 570 -521 580 -511
rect 1460 416 1468 425
rect 1478 416 1486 425
rect 1192 398 1200 405
rect 1214 395 1224 404
rect 1255 398 1263 406
rect 1278 397 1286 405
rect 1331 398 1339 406
rect 1351 396 1361 405
rect 1392 399 1400 407
rect 1415 398 1423 406
rect 233 -572 241 -563
rect 251 -572 259 -563
rect 300 -685 308 -678
rect 322 -688 332 -679
rect 363 -685 371 -677
rect 386 -686 394 -678
rect 426 -686 434 -678
rect 449 -687 457 -679
rect 494 -688 502 -680
rect 517 -689 525 -681
rect 565 -683 575 -673
rect 590 -682 600 -672
rect 232 -727 240 -718
rect 250 -727 258 -718
rect 309 -904 317 -897
rect 331 -907 341 -898
rect 372 -904 380 -896
rect 395 -905 403 -897
rect 435 -905 443 -897
rect 458 -906 466 -898
rect 503 -907 511 -899
rect 526 -908 534 -900
rect 562 -908 570 -900
rect 585 -909 593 -901
rect 635 -903 645 -893
rect 660 -902 670 -892
rect 1400 -421 1406 -416
rect 1419 -421 1426 -415
rect 1440 -421 1446 -416
rect 1459 -421 1466 -415
rect 1479 -422 1485 -416
rect 1498 -421 1505 -414
rect 1522 -422 1528 -416
rect 1540 -421 1547 -415
rect 1564 -421 1570 -416
rect 1582 -421 1589 -415
rect 232 -959 240 -950
rect 250 -959 258 -950
<< pdcontact >>
rect 375 1995 382 2001
rect 397 1991 406 1999
rect 441 1992 449 1999
rect 460 1991 468 1997
rect 545 1981 555 1991
rect 569 1978 579 1988
rect 285 1907 293 1916
rect 303 1907 312 1916
rect 1340 1906 1346 1912
rect 1359 1903 1365 1909
rect 1380 1903 1386 1909
rect 1400 1903 1406 1909
rect 1419 1903 1425 1909
rect 1438 1903 1444 1909
rect 1462 1903 1468 1909
rect 1481 1903 1487 1909
rect 1504 1906 1510 1912
rect 1522 1904 1529 1910
rect 375 1826 382 1832
rect 397 1822 406 1830
rect 441 1823 449 1830
rect 460 1822 468 1828
rect 504 1822 512 1829
rect 287 1745 295 1754
rect 305 1745 314 1754
rect 523 1821 531 1827
rect 600 1826 610 1836
rect 624 1823 634 1833
rect 355 1667 362 1673
rect 377 1663 386 1671
rect 421 1664 429 1671
rect 440 1663 448 1669
rect 484 1663 492 1670
rect 286 1590 294 1599
rect 304 1590 313 1599
rect 503 1662 511 1668
rect 552 1661 560 1668
rect 571 1660 579 1666
rect 620 1665 630 1675
rect 644 1662 654 1672
rect 364 1448 371 1454
rect 386 1444 395 1452
rect 430 1445 438 1452
rect 449 1444 457 1450
rect 493 1444 501 1451
rect 512 1443 520 1449
rect 561 1442 569 1449
rect 286 1358 294 1367
rect 304 1358 313 1367
rect 580 1441 588 1447
rect 620 1441 628 1448
rect 639 1440 647 1446
rect 690 1445 700 1455
rect 714 1442 724 1452
rect 244 1058 251 1064
rect 266 1054 275 1062
rect 310 1055 318 1062
rect 329 1054 337 1060
rect 447 1058 454 1064
rect 469 1054 478 1062
rect 513 1055 521 1062
rect 532 1054 540 1060
rect 634 1058 641 1064
rect 656 1054 665 1062
rect 700 1055 708 1062
rect 719 1054 727 1060
rect 815 1058 822 1064
rect 837 1054 846 1062
rect 881 1055 889 1062
rect 900 1054 908 1060
rect 971 1040 979 1049
rect 989 1040 998 1049
rect 250 769 257 775
rect 272 765 281 773
rect 316 766 324 773
rect 335 765 343 771
rect 453 769 460 775
rect 475 765 484 773
rect 519 766 527 773
rect 538 765 546 771
rect 640 769 647 775
rect 662 765 671 773
rect 706 766 714 773
rect 725 765 733 771
rect 821 769 828 775
rect 843 765 852 773
rect 887 766 895 773
rect 906 765 914 771
rect 973 748 981 757
rect 991 748 1000 757
rect 270 452 277 458
rect 292 448 301 456
rect 336 449 344 456
rect 355 448 363 454
rect 473 452 480 458
rect 495 448 504 456
rect 539 449 547 456
rect 558 448 566 454
rect 660 452 667 458
rect 682 448 691 456
rect 726 449 734 456
rect 745 448 753 454
rect 841 452 848 458
rect 863 448 872 456
rect 907 449 915 456
rect 926 448 934 454
rect 998 431 1006 440
rect 1016 431 1025 440
rect 268 161 275 167
rect 290 157 299 165
rect 334 158 342 165
rect 353 157 361 163
rect 471 161 478 167
rect 493 157 502 165
rect 537 158 545 165
rect 556 157 564 163
rect 658 161 665 167
rect 680 157 689 165
rect 724 158 732 165
rect 743 157 751 163
rect 839 161 846 167
rect 861 157 870 165
rect 905 158 913 165
rect 924 157 932 163
rect 1007 140 1015 149
rect 1025 140 1034 149
rect 321 -271 328 -265
rect 343 -275 352 -267
rect 387 -274 395 -267
rect 406 -275 414 -269
rect 491 -285 501 -275
rect 515 -288 525 -278
rect 231 -359 239 -350
rect 249 -359 258 -350
rect 321 -440 328 -434
rect 343 -444 352 -436
rect 387 -443 395 -436
rect 406 -444 414 -438
rect 450 -444 458 -437
rect 233 -521 241 -512
rect 251 -521 260 -512
rect 469 -445 477 -439
rect 546 -440 556 -430
rect 570 -443 580 -433
rect 1193 484 1200 490
rect 1215 480 1224 488
rect 1259 481 1267 488
rect 1278 480 1286 486
rect 1330 485 1337 491
rect 1352 481 1361 489
rect 1396 482 1404 489
rect 1415 481 1423 487
rect 1460 467 1468 476
rect 1478 467 1487 476
rect 301 -599 308 -593
rect 323 -603 332 -595
rect 367 -602 375 -595
rect 386 -603 394 -597
rect 430 -603 438 -596
rect 232 -676 240 -667
rect 250 -676 259 -667
rect 449 -604 457 -598
rect 498 -605 506 -598
rect 517 -606 525 -600
rect 566 -601 576 -591
rect 590 -604 600 -594
rect 310 -818 317 -812
rect 332 -822 341 -814
rect 376 -821 384 -814
rect 395 -822 403 -816
rect 439 -822 447 -815
rect 458 -823 466 -817
rect 507 -824 515 -817
rect 232 -908 240 -899
rect 250 -908 259 -899
rect 526 -825 534 -819
rect 566 -825 574 -818
rect 585 -826 593 -820
rect 636 -821 646 -811
rect 660 -824 670 -814
rect 1400 -360 1406 -354
rect 1419 -363 1425 -357
rect 1440 -363 1446 -357
rect 1460 -363 1466 -357
rect 1479 -363 1485 -357
rect 1498 -363 1504 -357
rect 1522 -363 1528 -357
rect 1541 -363 1547 -357
rect 1564 -360 1570 -354
rect 1582 -362 1589 -356
<< polysilicon >>
rect 386 2003 393 2006
rect 450 2003 457 2006
rect 559 1991 567 1997
rect 51 1956 295 1957
rect 386 1956 393 1988
rect 51 1944 393 1956
rect 51 1943 295 1944
rect 53 1927 67 1943
rect 53 258 66 1927
rect 295 1916 301 1919
rect 386 1918 393 1944
rect 450 1918 457 1988
rect 559 1944 567 1975
rect 525 1943 567 1944
rect 535 1934 567 1943
rect 295 1887 301 1907
rect 559 1913 567 1934
rect 1349 1914 1355 1918
rect 1390 1914 1396 1918
rect 1429 1914 1435 1918
rect 1472 1914 1478 1918
rect 1514 1914 1520 1918
rect 386 1899 393 1903
rect 300 1880 301 1887
rect 295 1865 301 1880
rect 450 1888 457 1903
rect 559 1889 567 1897
rect 1349 1892 1355 1903
rect 295 1853 301 1856
rect 1349 1853 1355 1886
rect 1390 1853 1396 1903
rect 1429 1853 1435 1903
rect 1472 1853 1478 1903
rect 1514 1881 1520 1903
rect 1500 1875 1520 1881
rect 1514 1853 1520 1875
rect 386 1834 393 1837
rect 450 1834 457 1837
rect 614 1836 622 1842
rect 1349 1837 1355 1842
rect 513 1833 520 1836
rect 80 1787 356 1788
rect 386 1787 393 1819
rect 80 1775 393 1787
rect 81 1616 94 1775
rect 297 1754 303 1757
rect 386 1749 393 1775
rect 450 1749 457 1819
rect 297 1725 303 1745
rect 513 1748 520 1818
rect 614 1789 622 1820
rect 580 1788 622 1789
rect 590 1779 622 1788
rect 1390 1792 1396 1842
rect 614 1758 622 1779
rect 386 1730 393 1734
rect 302 1718 303 1725
rect 297 1703 303 1718
rect 450 1719 457 1734
rect 614 1734 622 1742
rect 513 1715 520 1733
rect 1068 1715 1083 1718
rect 512 1705 1083 1715
rect 297 1691 303 1694
rect 366 1675 373 1678
rect 430 1675 437 1678
rect 493 1674 500 1677
rect 634 1675 642 1681
rect 366 1632 373 1660
rect 108 1616 373 1632
rect 82 528 92 1616
rect 108 1609 121 1616
rect 108 846 120 1609
rect 296 1599 302 1602
rect 366 1590 373 1616
rect 430 1590 437 1660
rect 561 1672 568 1675
rect 296 1570 302 1590
rect 493 1589 500 1659
rect 366 1571 373 1575
rect 301 1563 302 1570
rect 296 1548 302 1563
rect 430 1560 437 1575
rect 561 1587 568 1657
rect 634 1628 642 1659
rect 600 1627 642 1628
rect 610 1618 642 1627
rect 634 1597 642 1618
rect 493 1556 500 1574
rect 634 1573 642 1581
rect 520 1556 530 1557
rect 492 1546 530 1556
rect 561 1554 568 1572
rect 296 1536 302 1539
rect 520 1535 530 1546
rect 560 1544 581 1554
rect 596 1544 597 1554
rect 1068 1535 1083 1705
rect 1429 1628 1435 1842
rect 1429 1612 1435 1621
rect 520 1522 1083 1535
rect 375 1456 382 1459
rect 439 1456 446 1459
rect 502 1455 509 1458
rect 337 1410 342 1412
rect 190 1397 221 1410
rect 234 1409 355 1410
rect 375 1409 382 1441
rect 234 1397 382 1409
rect 190 1131 199 1397
rect 375 1371 382 1397
rect 439 1371 446 1441
rect 570 1453 577 1456
rect 296 1367 302 1370
rect 296 1338 302 1358
rect 502 1370 509 1440
rect 629 1452 636 1493
rect 704 1455 712 1461
rect 375 1352 382 1356
rect 301 1331 302 1338
rect 296 1316 302 1331
rect 439 1341 446 1356
rect 570 1368 577 1438
rect 502 1337 509 1355
rect 629 1367 636 1437
rect 704 1408 712 1439
rect 670 1407 712 1408
rect 680 1398 712 1407
rect 704 1377 712 1398
rect 529 1337 539 1338
rect 501 1327 539 1337
rect 570 1335 577 1353
rect 704 1353 712 1361
rect 629 1346 636 1352
rect 529 1316 539 1327
rect 569 1325 590 1335
rect 605 1325 606 1335
rect 1068 1316 1083 1522
rect 1097 1556 1111 1564
rect 1097 1545 1098 1556
rect 1097 1337 1111 1545
rect 1126 1506 1140 1509
rect 296 1304 302 1307
rect 529 1303 1086 1316
rect 190 1123 666 1131
rect 190 1120 326 1123
rect 190 1119 199 1120
rect 188 1095 205 1103
rect 215 1095 216 1103
rect 188 1092 216 1095
rect 206 1016 216 1092
rect 255 1066 262 1069
rect 319 1066 326 1120
rect 458 1066 465 1069
rect 522 1066 529 1069
rect 645 1066 652 1123
rect 709 1066 716 1069
rect 826 1066 833 1099
rect 890 1066 897 1069
rect 255 1016 262 1051
rect 206 1008 262 1016
rect 206 1007 216 1008
rect 255 981 262 1008
rect 319 981 326 1051
rect 458 981 465 1051
rect 522 981 529 1051
rect 645 981 652 1051
rect 709 981 716 1051
rect 826 981 833 1051
rect 890 981 897 1051
rect 981 1049 987 1052
rect 981 1024 987 1040
rect 986 1015 987 1024
rect 981 998 987 1015
rect 981 986 987 989
rect 255 922 262 966
rect 319 961 326 966
rect 458 922 465 966
rect 522 937 529 966
rect 645 962 652 966
rect 709 938 716 966
rect 826 962 833 966
rect 255 915 465 922
rect 890 919 897 966
rect 121 834 672 842
rect 121 831 332 834
rect 204 803 222 814
rect 212 727 222 803
rect 261 777 268 780
rect 325 777 332 831
rect 464 777 471 780
rect 528 777 535 780
rect 651 777 658 834
rect 715 777 722 780
rect 832 777 839 810
rect 896 777 903 780
rect 261 727 268 762
rect 212 719 268 727
rect 212 718 222 719
rect 261 692 268 719
rect 325 692 332 762
rect 464 692 471 762
rect 528 692 535 762
rect 651 692 658 762
rect 715 692 722 762
rect 832 692 839 762
rect 896 692 903 762
rect 983 757 989 760
rect 983 732 989 748
rect 988 723 989 732
rect 983 706 989 723
rect 983 694 989 697
rect 261 633 268 677
rect 325 672 332 677
rect 464 633 471 677
rect 528 648 535 677
rect 651 673 658 677
rect 715 649 722 677
rect 832 673 839 677
rect 261 626 471 633
rect 896 630 903 677
rect 92 525 223 526
rect 92 517 692 525
rect 92 514 352 517
rect 226 487 242 497
rect 214 486 242 487
rect 232 410 242 486
rect 281 460 288 463
rect 345 460 352 514
rect 484 460 491 463
rect 548 460 555 463
rect 671 460 678 517
rect 735 460 742 463
rect 852 460 859 493
rect 916 460 923 463
rect 281 410 288 445
rect 232 402 288 410
rect 232 401 242 402
rect 281 375 288 402
rect 345 375 352 445
rect 484 375 491 445
rect 548 375 555 445
rect 671 375 678 445
rect 735 375 742 445
rect 852 375 859 445
rect 916 375 923 445
rect 1008 440 1014 443
rect 1008 415 1014 431
rect 1013 406 1014 415
rect 1008 389 1014 406
rect 1008 377 1014 380
rect 281 316 288 360
rect 345 355 352 360
rect 484 316 491 360
rect 548 331 555 360
rect 671 356 678 360
rect 735 332 742 360
rect 852 356 859 360
rect 281 309 491 316
rect 916 313 923 360
rect 51 234 66 258
rect 51 226 690 234
rect 51 223 350 226
rect 51 222 66 223
rect 51 0 65 222
rect 107 0 108 18
rect 107 -585 118 0
rect 162 -379 176 223
rect 212 205 240 206
rect 212 195 215 205
rect 228 195 240 205
rect 230 122 240 195
rect 279 169 286 172
rect 343 169 350 223
rect 482 169 489 172
rect 546 169 553 172
rect 669 169 676 226
rect 733 169 740 172
rect 850 169 857 202
rect 914 169 921 172
rect 230 119 254 122
rect 279 119 286 154
rect 230 111 286 119
rect 230 110 254 111
rect 239 0 254 110
rect 279 84 286 111
rect 343 84 350 154
rect 482 84 489 154
rect 546 84 553 154
rect 669 84 676 154
rect 733 84 740 154
rect 850 84 857 154
rect 914 84 921 154
rect 1017 149 1023 152
rect 1017 124 1023 140
rect 1022 115 1023 124
rect 1017 98 1023 115
rect 1068 124 1083 1303
rect 1097 415 1111 1325
rect 1110 406 1111 415
rect 1068 115 1069 124
rect 1017 86 1023 89
rect 279 25 286 69
rect 343 64 350 69
rect 482 25 489 69
rect 546 40 553 69
rect 669 65 676 69
rect 733 41 740 69
rect 850 65 857 69
rect 279 18 489 25
rect 914 22 921 69
rect 332 -263 339 -260
rect 396 -263 403 -260
rect 505 -275 513 -269
rect 216 -309 222 -308
rect 216 -310 241 -309
rect 332 -310 339 -278
rect 242 -322 339 -310
rect 216 -323 241 -322
rect 216 -324 222 -323
rect 241 -350 247 -347
rect 332 -348 339 -322
rect 396 -348 403 -278
rect 505 -322 513 -291
rect 471 -323 513 -322
rect 481 -332 513 -323
rect 241 -379 247 -359
rect 505 -353 513 -332
rect 332 -367 339 -363
rect 162 -386 216 -379
rect 246 -386 247 -379
rect 241 -401 247 -386
rect 396 -378 403 -363
rect 505 -377 513 -369
rect 241 -413 247 -410
rect 332 -432 339 -429
rect 396 -432 403 -429
rect 560 -430 568 -424
rect 459 -433 466 -430
rect 217 -479 302 -478
rect 332 -479 339 -447
rect 217 -491 339 -479
rect 243 -512 249 -509
rect 332 -517 339 -491
rect 396 -517 403 -447
rect 243 -541 249 -521
rect 459 -518 466 -448
rect 560 -477 568 -446
rect 526 -478 568 -477
rect 536 -487 568 -478
rect 560 -508 568 -487
rect 332 -536 339 -532
rect 248 -548 249 -541
rect 243 -563 249 -548
rect 396 -547 403 -532
rect 560 -532 568 -524
rect 459 -551 466 -533
rect 1068 -548 1083 115
rect 1097 15 1111 406
rect 1126 509 1140 1493
rect 1472 1411 1478 1842
rect 1514 1837 1520 1842
rect 1341 1024 1347 1043
rect 1126 501 1127 509
rect 1126 25 1140 501
rect 1341 603 1347 1015
rect 1204 492 1211 495
rect 1268 492 1275 495
rect 1341 493 1348 603
rect 1405 493 1412 496
rect 1204 436 1211 477
rect 1210 427 1211 436
rect 1204 407 1211 427
rect 1268 407 1275 477
rect 1341 408 1348 478
rect 1405 408 1412 478
rect 1470 476 1476 479
rect 1470 447 1476 467
rect 1475 437 1476 447
rect 1470 425 1476 437
rect 1470 413 1476 416
rect 1204 388 1211 392
rect 1268 319 1275 392
rect 1341 389 1348 393
rect 1405 390 1412 393
rect 1405 338 1413 390
rect 1412 327 1413 338
rect 1269 123 1275 319
rect 1269 91 1275 116
rect 1068 -551 1084 -548
rect 458 -561 1084 -551
rect 1068 -562 1084 -561
rect 243 -575 249 -572
rect 107 -695 119 -585
rect 312 -591 319 -588
rect 376 -591 383 -588
rect 439 -592 446 -589
rect 580 -591 588 -585
rect 312 -634 319 -606
rect 217 -650 319 -634
rect 242 -667 248 -664
rect 312 -676 319 -650
rect 376 -676 383 -606
rect 507 -594 514 -591
rect 107 -702 197 -695
rect 107 -703 211 -702
rect 242 -696 248 -676
rect 439 -677 446 -607
rect 312 -695 319 -691
rect 247 -703 248 -696
rect 107 -708 119 -703
rect 242 -718 248 -703
rect 376 -706 383 -691
rect 507 -679 514 -609
rect 580 -638 588 -607
rect 546 -639 588 -638
rect 556 -648 588 -639
rect 580 -669 588 -648
rect 439 -710 446 -692
rect 580 -693 588 -685
rect 466 -710 476 -709
rect 438 -720 476 -710
rect 507 -712 514 -694
rect 242 -730 248 -727
rect 466 -731 476 -720
rect 506 -722 527 -712
rect 542 -722 543 -712
rect 1069 -731 1084 -562
rect 466 -744 1084 -731
rect 1096 -710 1112 15
rect 1096 -721 1099 -710
rect 1096 -735 1112 -721
rect 321 -810 328 -807
rect 385 -810 392 -807
rect 448 -811 455 -808
rect 283 -856 288 -854
rect 211 -857 301 -856
rect 321 -857 328 -825
rect 211 -869 328 -857
rect 321 -895 328 -869
rect 385 -895 392 -825
rect 516 -813 523 -810
rect 242 -899 248 -896
rect 242 -928 248 -908
rect 448 -896 455 -826
rect 575 -814 582 -773
rect 650 -811 658 -805
rect 321 -914 328 -910
rect 247 -935 248 -928
rect 242 -950 248 -935
rect 385 -925 392 -910
rect 516 -898 523 -828
rect 448 -929 455 -911
rect 575 -899 582 -829
rect 650 -858 658 -827
rect 616 -859 658 -858
rect 626 -868 658 -859
rect 650 -889 658 -868
rect 475 -929 485 -928
rect 447 -939 485 -929
rect 516 -931 523 -913
rect 650 -913 658 -905
rect 575 -920 582 -914
rect 475 -950 485 -939
rect 515 -941 536 -931
rect 551 -941 552 -931
rect 1069 -950 1084 -744
rect 1098 -929 1112 -735
rect 1126 -760 1141 25
rect 1409 -352 1415 -348
rect 1450 -352 1456 -348
rect 1489 -352 1495 -348
rect 1532 -352 1538 -348
rect 1574 -352 1580 -348
rect 1409 -374 1415 -363
rect 1409 -413 1415 -380
rect 1450 -413 1456 -363
rect 1489 -413 1495 -363
rect 1532 -413 1538 -363
rect 1574 -385 1580 -363
rect 1560 -391 1580 -385
rect 1574 -413 1580 -391
rect 1409 -429 1415 -424
rect 1450 -474 1456 -424
rect 1489 -638 1495 -424
rect 1489 -654 1495 -645
rect 1126 -773 1127 -760
rect 1126 -792 1141 -773
rect 242 -962 248 -959
rect 475 -963 1087 -950
rect 1069 -1001 1084 -963
rect 1098 -1001 1112 -941
rect 1127 -1001 1141 -792
rect 1532 -855 1538 -424
rect 1574 -429 1580 -424
<< polycontact >>
rect 524 1933 535 1943
rect 295 1880 300 1887
rect 450 1876 458 1888
rect 1349 1886 1355 1892
rect 1495 1875 1500 1881
rect 579 1778 590 1788
rect 1390 1781 1397 1792
rect 297 1718 302 1725
rect 450 1707 458 1719
rect 296 1563 301 1570
rect 599 1617 610 1627
rect 430 1548 438 1560
rect 581 1543 596 1554
rect 1428 1621 1435 1628
rect 628 1493 637 1503
rect 221 1397 234 1410
rect 296 1331 301 1338
rect 439 1329 447 1341
rect 669 1397 680 1407
rect 590 1324 605 1335
rect 1098 1545 1113 1556
rect 1126 1493 1142 1506
rect 1096 1325 1113 1337
rect 205 1095 215 1103
rect 826 1099 833 1106
rect 981 1015 986 1024
rect 522 929 529 937
rect 709 930 716 938
rect 890 912 897 919
rect 107 830 121 846
rect 194 803 204 814
rect 832 810 839 817
rect 983 723 988 732
rect 528 640 535 648
rect 715 641 722 649
rect 896 623 903 630
rect 82 513 92 528
rect 213 487 226 497
rect 852 493 859 500
rect 1008 406 1013 415
rect 548 323 555 331
rect 735 324 742 332
rect 916 306 923 313
rect 108 0 118 18
rect 215 195 228 205
rect 850 202 857 209
rect 1017 115 1022 124
rect 1096 406 1110 415
rect 1069 115 1083 124
rect 546 32 553 40
rect 733 33 740 41
rect 914 15 921 22
rect 216 -322 242 -310
rect 470 -333 481 -323
rect 216 -386 225 -379
rect 241 -386 246 -379
rect 396 -390 404 -378
rect 197 -491 217 -478
rect 525 -488 536 -478
rect 243 -548 248 -541
rect 396 -559 404 -547
rect 1472 1400 1478 1411
rect 1340 1015 1348 1024
rect 1127 501 1140 509
rect 1204 427 1210 436
rect 1470 437 1475 447
rect 1405 327 1412 338
rect 1268 116 1276 123
rect 197 -650 217 -634
rect 197 -702 211 -695
rect 242 -703 247 -696
rect 545 -649 556 -639
rect 376 -718 384 -706
rect 527 -723 542 -712
rect 1099 -721 1114 -710
rect 574 -773 583 -763
rect 197 -869 211 -856
rect 242 -935 247 -928
rect 385 -937 393 -925
rect 615 -869 626 -859
rect 536 -942 551 -931
rect 1409 -380 1415 -374
rect 1555 -391 1560 -385
rect 1450 -485 1457 -474
rect 1488 -645 1495 -638
rect 1127 -773 1143 -760
rect 1097 -941 1114 -929
rect 1532 -866 1538 -855
<< metal1 >>
rect 441 2021 449 2026
rect 375 2015 449 2021
rect 375 2001 382 2015
rect 441 1999 449 2015
rect 581 2011 589 2019
rect 546 2005 589 2011
rect 397 1960 406 1991
rect 546 1991 554 2005
rect 460 1960 468 1991
rect 397 1958 468 1960
rect 397 1957 469 1958
rect 397 1952 494 1957
rect 460 1948 494 1952
rect 286 1916 293 1932
rect 396 1924 445 1932
rect 133 1887 142 1895
rect 303 1887 311 1907
rect 374 1890 382 1909
rect 396 1915 406 1924
rect 437 1917 445 1924
rect 460 1916 468 1948
rect 483 1943 494 1948
rect 569 1945 579 1978
rect 588 1945 1100 1946
rect 483 1933 524 1943
rect 569 1936 1100 1945
rect 569 1910 579 1936
rect 588 1935 1100 1936
rect 133 1880 295 1887
rect 133 1868 142 1880
rect 235 1879 273 1880
rect 131 1799 142 1868
rect 303 1876 450 1887
rect 545 1883 554 1899
rect 1092 1893 1100 1935
rect 1340 1922 1363 1928
rect 1340 1912 1346 1922
rect 1504 1912 1510 1928
rect 1092 1892 1356 1893
rect 1092 1886 1349 1892
rect 1355 1886 1356 1892
rect 1359 1890 1365 1903
rect 1380 1890 1386 1903
rect 1359 1884 1386 1890
rect 1400 1890 1406 1903
rect 1419 1890 1425 1903
rect 1400 1884 1425 1890
rect 1438 1890 1444 1903
rect 1462 1890 1468 1903
rect 1438 1884 1468 1890
rect 545 1877 580 1883
rect 1481 1881 1487 1903
rect 1522 1882 1529 1904
rect 1522 1881 1536 1882
rect 1609 1881 1674 1882
rect 303 1875 458 1876
rect 1481 1875 1495 1881
rect 1522 1876 1674 1881
rect 303 1865 311 1875
rect 1481 1869 1487 1875
rect 286 1846 293 1856
rect 441 1852 449 1857
rect 636 1856 644 1864
rect 375 1851 499 1852
rect 504 1851 512 1856
rect 375 1846 512 1851
rect 375 1832 382 1846
rect 441 1845 512 1846
rect 441 1830 449 1845
rect 504 1829 512 1845
rect 601 1850 644 1856
rect 1359 1863 1487 1869
rect 1359 1851 1366 1863
rect 601 1836 609 1850
rect 1399 1851 1406 1863
rect 1438 1852 1445 1863
rect 131 1772 141 1799
rect 397 1791 406 1822
rect 460 1791 468 1822
rect 397 1790 468 1791
rect 523 1790 531 1821
rect 397 1788 531 1790
rect 1340 1831 1346 1845
rect 1380 1831 1386 1845
rect 1480 1851 1487 1863
rect 1419 1831 1425 1844
rect 1522 1851 1529 1876
rect 1462 1831 1468 1844
rect 1340 1826 1468 1831
rect 1504 1828 1510 1845
rect 624 1790 634 1823
rect 639 1790 1390 1791
rect 397 1787 532 1788
rect 572 1787 579 1788
rect 397 1783 579 1787
rect 460 1779 579 1783
rect 523 1778 579 1779
rect 624 1781 1390 1790
rect 131 1769 142 1772
rect 11 1231 35 1232
rect 0 1218 40 1231
rect 0 -855 9 1218
rect 108 846 120 847
rect 82 70 92 513
rect 82 -541 93 70
rect 108 18 120 830
rect 133 205 142 1769
rect 288 1754 295 1769
rect 396 1755 445 1763
rect 155 1718 297 1725
rect 305 1718 313 1745
rect 374 1722 382 1740
rect 396 1746 406 1755
rect 437 1748 445 1755
rect 460 1754 508 1762
rect 460 1747 468 1754
rect 500 1747 508 1754
rect 523 1746 531 1778
rect 624 1755 634 1781
rect 600 1728 609 1744
rect 600 1722 635 1728
rect 155 497 163 1718
rect 235 1717 270 1718
rect 305 1707 450 1718
rect 305 1706 458 1707
rect 305 1703 313 1706
rect 288 1684 295 1694
rect 421 1693 429 1698
rect 355 1692 479 1693
rect 484 1692 492 1697
rect 656 1695 664 1703
rect 355 1691 492 1692
rect 355 1690 547 1691
rect 552 1690 560 1695
rect 355 1687 560 1690
rect 355 1673 362 1687
rect 421 1686 560 1687
rect 421 1671 429 1686
rect 484 1684 560 1686
rect 484 1670 492 1684
rect 377 1632 386 1663
rect 552 1668 560 1684
rect 621 1689 664 1695
rect 621 1675 629 1689
rect 440 1632 448 1663
rect 377 1631 448 1632
rect 503 1631 511 1662
rect 377 1629 511 1631
rect 571 1629 579 1660
rect 377 1628 512 1629
rect 527 1628 579 1629
rect 377 1627 579 1628
rect 644 1629 654 1662
rect 644 1628 1437 1629
rect 377 1626 580 1627
rect 592 1626 599 1627
rect 377 1624 599 1626
rect 440 1620 599 1624
rect 503 1619 599 1620
rect 535 1618 599 1619
rect 571 1617 599 1618
rect 644 1621 1428 1628
rect 1435 1621 1437 1628
rect 644 1620 671 1621
rect 287 1599 294 1615
rect 376 1596 425 1604
rect 233 1570 268 1571
rect 174 1563 296 1570
rect 304 1568 312 1590
rect 174 816 182 1563
rect 304 1559 336 1568
rect 354 1563 362 1581
rect 376 1587 386 1596
rect 417 1589 425 1596
rect 440 1595 488 1603
rect 503 1601 511 1602
rect 440 1588 448 1595
rect 480 1588 488 1595
rect 502 1594 556 1601
rect 503 1587 511 1594
rect 535 1593 556 1594
rect 548 1586 556 1593
rect 571 1585 579 1617
rect 644 1594 654 1620
rect 620 1567 629 1583
rect 620 1561 655 1567
rect 304 1558 430 1559
rect 304 1548 312 1558
rect 328 1548 430 1558
rect 974 1556 1114 1557
rect 974 1554 1098 1556
rect 329 1547 438 1548
rect 596 1545 1098 1554
rect 1113 1545 1114 1556
rect 596 1544 1114 1545
rect 287 1529 294 1539
rect 626 1503 1126 1505
rect 626 1493 628 1503
rect 637 1493 1126 1503
rect 626 1492 1141 1493
rect 430 1474 438 1479
rect 364 1473 488 1474
rect 493 1473 501 1478
rect 364 1472 501 1473
rect 364 1471 556 1472
rect 561 1471 569 1476
rect 726 1475 734 1483
rect 620 1471 628 1475
rect 364 1468 628 1471
rect 364 1454 371 1468
rect 430 1467 628 1468
rect 430 1452 438 1467
rect 493 1465 628 1467
rect 493 1451 501 1465
rect 559 1464 628 1465
rect 221 1410 233 1421
rect 386 1413 395 1444
rect 561 1449 569 1464
rect 449 1413 457 1444
rect 386 1412 457 1413
rect 512 1412 520 1443
rect 620 1448 628 1464
rect 691 1469 734 1475
rect 691 1455 699 1469
rect 386 1410 520 1412
rect 580 1410 588 1441
rect 386 1409 521 1410
rect 536 1409 588 1410
rect 639 1409 647 1440
rect 386 1407 647 1409
rect 714 1409 724 1442
rect 728 1409 1472 1411
rect 386 1406 648 1407
rect 660 1406 669 1407
rect 386 1405 669 1406
rect 449 1401 669 1405
rect 512 1400 669 1401
rect 544 1399 669 1400
rect 580 1398 669 1399
rect 639 1397 669 1398
rect 714 1401 1472 1409
rect 714 1400 741 1401
rect 1478 1401 1531 1411
rect 287 1367 294 1383
rect 385 1377 434 1385
rect 304 1341 312 1358
rect 337 1341 345 1342
rect 363 1341 371 1362
rect 385 1368 395 1377
rect 426 1370 434 1377
rect 449 1376 497 1384
rect 512 1382 520 1383
rect 449 1369 457 1376
rect 489 1369 497 1376
rect 511 1375 565 1382
rect 512 1368 520 1375
rect 544 1374 565 1375
rect 557 1367 565 1374
rect 580 1380 588 1381
rect 603 1380 624 1381
rect 580 1373 624 1380
rect 580 1366 588 1373
rect 616 1366 624 1373
rect 639 1365 647 1397
rect 714 1374 724 1400
rect 690 1347 699 1363
rect 690 1341 725 1347
rect 304 1340 389 1341
rect 228 1338 270 1339
rect 203 1331 296 1338
rect 205 1231 215 1331
rect 304 1330 439 1340
rect 304 1316 312 1330
rect 337 1329 439 1330
rect 900 1337 1112 1338
rect 900 1336 1096 1337
rect 685 1335 1096 1336
rect 338 1328 447 1329
rect 605 1325 1096 1335
rect 287 1297 294 1307
rect 214 1218 215 1231
rect 205 1103 215 1218
rect 575 1106 834 1108
rect 261 1095 560 1105
rect 575 1099 826 1106
rect 833 1099 834 1106
rect 575 1098 834 1099
rect 310 1084 318 1095
rect 513 1084 521 1095
rect 244 1078 318 1084
rect 244 1064 251 1078
rect 310 1062 318 1078
rect 447 1078 521 1084
rect 447 1064 454 1078
rect 266 1023 275 1054
rect 513 1062 521 1078
rect 329 1033 337 1054
rect 328 1023 337 1033
rect 266 1020 337 1023
rect 469 1023 478 1054
rect 532 1023 540 1054
rect 469 1022 540 1023
rect 576 1022 585 1098
rect 700 1084 708 1093
rect 881 1084 889 1093
rect 634 1078 708 1084
rect 634 1064 641 1078
rect 700 1062 708 1078
rect 266 1015 363 1020
rect 469 1015 585 1022
rect 815 1078 889 1084
rect 815 1064 822 1078
rect 656 1023 665 1054
rect 881 1062 889 1078
rect 719 1023 727 1054
rect 656 1022 727 1023
rect 837 1023 846 1054
rect 900 1023 908 1054
rect 972 1049 979 1065
rect 989 1024 997 1040
rect 837 1022 908 1023
rect 914 1022 981 1024
rect 656 1015 773 1022
rect 837 1015 981 1022
rect 989 1015 1340 1024
rect 329 1011 363 1015
rect 265 987 314 995
rect 243 950 251 972
rect 265 978 275 987
rect 306 980 314 987
rect 329 979 337 1011
rect 352 938 363 1011
rect 532 1013 585 1015
rect 719 1013 773 1015
rect 468 987 517 995
rect 446 950 454 972
rect 468 978 478 987
rect 509 980 517 987
rect 532 979 540 1013
rect 655 987 704 995
rect 633 950 641 972
rect 655 978 665 987
rect 696 980 704 987
rect 719 979 727 1013
rect 352 937 709 938
rect 352 929 522 937
rect 529 930 709 937
rect 716 930 750 938
rect 529 929 750 930
rect 352 927 750 929
rect 761 919 773 1013
rect 900 1013 928 1015
rect 836 987 885 995
rect 814 950 822 972
rect 836 978 846 987
rect 877 980 885 987
rect 900 979 908 1013
rect 989 998 997 1015
rect 972 979 979 989
rect 761 912 890 919
rect 897 912 930 919
rect 761 909 930 912
rect 581 817 840 819
rect 184 803 194 814
rect 267 806 566 816
rect 581 810 832 817
rect 839 810 840 817
rect 581 809 840 810
rect 316 795 324 806
rect 519 795 527 806
rect 250 789 324 795
rect 250 775 257 789
rect 316 773 324 789
rect 453 789 527 795
rect 453 775 460 789
rect 272 734 281 765
rect 519 773 527 789
rect 335 744 343 765
rect 334 734 343 744
rect 272 731 343 734
rect 475 734 484 765
rect 538 734 546 765
rect 475 733 546 734
rect 582 733 591 809
rect 706 795 714 804
rect 887 795 895 804
rect 640 789 714 795
rect 640 775 647 789
rect 706 773 714 789
rect 272 726 369 731
rect 475 726 591 733
rect 821 789 895 795
rect 821 775 828 789
rect 662 734 671 765
rect 887 773 895 789
rect 725 734 733 765
rect 662 733 733 734
rect 843 734 852 765
rect 906 734 914 765
rect 974 757 981 773
rect 843 733 914 734
rect 932 733 961 734
rect 662 726 779 733
rect 843 732 961 733
rect 991 732 999 748
rect 843 726 983 732
rect 335 722 369 726
rect 271 698 320 706
rect 249 661 257 683
rect 271 689 281 698
rect 312 691 320 698
rect 335 690 343 722
rect 358 649 369 722
rect 538 724 591 726
rect 725 724 779 726
rect 474 698 523 706
rect 452 661 460 683
rect 474 689 484 698
rect 515 691 523 698
rect 538 690 546 724
rect 661 698 710 706
rect 639 661 647 683
rect 661 689 671 698
rect 702 691 710 698
rect 725 690 733 724
rect 358 648 715 649
rect 358 640 528 648
rect 535 641 715 648
rect 722 641 756 649
rect 535 640 756 641
rect 358 638 756 640
rect 767 630 779 724
rect 906 724 983 726
rect 842 698 891 706
rect 820 661 828 683
rect 842 689 852 698
rect 883 691 891 698
rect 906 690 914 724
rect 932 723 983 724
rect 991 723 1024 732
rect 991 706 999 723
rect 974 687 981 697
rect 1011 648 1022 723
rect 767 623 896 630
rect 903 623 936 630
rect 767 620 936 623
rect 1012 509 1021 648
rect 1259 511 1267 515
rect 1396 511 1404 516
rect 1259 510 1404 511
rect 601 500 860 502
rect 1012 501 1127 509
rect 1140 501 1142 509
rect 155 495 213 497
rect 161 488 213 495
rect 155 487 213 488
rect 287 489 586 499
rect 601 493 852 500
rect 859 493 860 500
rect 601 492 860 493
rect 336 478 344 489
rect 539 478 547 489
rect 270 472 344 478
rect 270 458 277 472
rect 336 456 344 472
rect 473 472 547 478
rect 473 458 480 472
rect 292 417 301 448
rect 539 456 547 472
rect 355 427 363 448
rect 354 417 363 427
rect 292 414 363 417
rect 495 417 504 448
rect 558 417 566 448
rect 495 416 566 417
rect 602 416 611 492
rect 726 478 734 487
rect 907 478 915 487
rect 660 472 734 478
rect 660 458 667 472
rect 726 456 734 472
rect 292 409 389 414
rect 495 409 611 416
rect 841 472 915 478
rect 841 458 848 472
rect 682 417 691 448
rect 907 456 915 472
rect 745 417 753 448
rect 682 416 753 417
rect 863 417 872 448
rect 926 417 934 448
rect 999 440 1006 456
rect 1135 436 1142 501
rect 1193 506 1404 510
rect 1193 504 1267 506
rect 1193 490 1200 504
rect 1259 488 1267 504
rect 1330 505 1404 506
rect 1330 491 1337 505
rect 1215 449 1224 480
rect 1396 489 1404 505
rect 1278 449 1286 480
rect 1215 447 1286 449
rect 1352 450 1361 481
rect 1415 450 1423 481
rect 1461 476 1468 492
rect 1352 448 1423 450
rect 1478 449 1486 467
rect 1352 447 1424 448
rect 1215 446 1287 447
rect 1297 446 1470 447
rect 1215 442 1470 446
rect 1215 441 1361 442
rect 1278 440 1361 441
rect 1278 438 1299 440
rect 1415 438 1470 442
rect 863 416 934 417
rect 682 409 799 416
rect 863 415 969 416
rect 1016 415 1024 431
rect 1135 427 1204 436
rect 1210 427 1213 436
rect 1068 415 1142 416
rect 863 409 1008 415
rect 355 405 389 409
rect 291 381 340 389
rect 269 344 277 366
rect 291 372 301 381
rect 332 374 340 381
rect 355 373 363 405
rect 378 332 389 405
rect 558 407 611 409
rect 745 407 799 409
rect 494 381 543 389
rect 472 344 480 366
rect 494 372 504 381
rect 535 374 543 381
rect 558 373 566 407
rect 681 381 730 389
rect 659 344 667 366
rect 681 372 691 381
rect 722 374 730 381
rect 745 373 753 407
rect 378 331 735 332
rect 378 323 548 331
rect 555 324 735 331
rect 742 324 776 332
rect 555 323 776 324
rect 378 321 776 323
rect 787 313 799 407
rect 926 407 1008 409
rect 862 381 911 389
rect 840 344 848 366
rect 862 372 872 381
rect 903 374 911 381
rect 926 373 934 407
rect 943 406 1008 407
rect 1016 406 1096 415
rect 1110 406 1142 415
rect 1016 389 1024 406
rect 999 370 1006 380
rect 1135 338 1142 406
rect 1214 413 1263 421
rect 1192 376 1200 398
rect 1214 404 1224 413
rect 1255 406 1263 413
rect 1278 415 1339 424
rect 1278 405 1286 415
rect 1331 406 1339 415
rect 1351 414 1400 422
rect 1351 405 1361 414
rect 1392 407 1400 414
rect 1415 406 1423 438
rect 1431 437 1470 438
rect 1478 439 1674 449
rect 1478 425 1486 439
rect 1461 406 1468 416
rect 1135 327 1405 338
rect 1412 327 1415 338
rect 787 306 916 313
rect 923 306 956 313
rect 787 303 956 306
rect 599 209 858 211
rect 133 195 215 205
rect 285 198 584 208
rect 599 202 850 209
rect 857 202 858 209
rect 599 201 858 202
rect 118 0 120 18
rect 191 -309 201 195
rect 334 187 342 198
rect 537 187 545 198
rect 268 181 342 187
rect 268 167 275 181
rect 334 165 342 181
rect 471 181 545 187
rect 471 167 478 181
rect 290 126 299 157
rect 537 165 545 181
rect 353 136 361 157
rect 352 126 361 136
rect 290 123 361 126
rect 493 126 502 157
rect 556 126 564 157
rect 493 125 564 126
rect 600 125 609 201
rect 724 187 732 196
rect 905 187 913 196
rect 658 181 732 187
rect 658 167 665 181
rect 724 165 732 181
rect 290 118 387 123
rect 493 118 609 125
rect 839 181 913 187
rect 839 167 846 181
rect 680 126 689 157
rect 905 165 913 181
rect 743 126 751 157
rect 680 125 751 126
rect 861 126 870 157
rect 924 126 932 157
rect 1008 149 1015 165
rect 861 125 932 126
rect 680 118 797 125
rect 861 124 952 125
rect 1025 124 1033 140
rect 1068 124 1085 125
rect 861 118 1017 124
rect 353 114 387 118
rect 289 90 338 98
rect 267 53 275 75
rect 289 81 299 90
rect 330 83 338 90
rect 353 82 361 114
rect 376 41 387 114
rect 556 116 609 118
rect 743 116 797 118
rect 492 90 541 98
rect 470 53 478 75
rect 492 81 502 90
rect 533 83 541 90
rect 556 82 564 116
rect 679 90 728 98
rect 657 53 665 75
rect 679 81 689 90
rect 720 83 728 90
rect 743 82 751 116
rect 376 40 733 41
rect 376 32 546 40
rect 553 33 733 40
rect 740 33 774 41
rect 553 32 774 33
rect 376 30 774 32
rect 785 22 797 116
rect 924 116 1017 118
rect 860 90 909 98
rect 838 53 846 75
rect 860 81 870 90
rect 901 83 909 90
rect 924 82 932 116
rect 986 115 1017 116
rect 1025 115 1069 124
rect 1083 123 1276 124
rect 1083 116 1268 123
rect 1083 115 1085 116
rect 1025 98 1033 115
rect 1008 79 1015 89
rect 785 15 914 22
rect 921 15 954 22
rect 785 12 954 15
rect 387 -245 395 -240
rect 321 -251 395 -245
rect 321 -265 328 -251
rect 387 -267 395 -251
rect 527 -255 535 -247
rect 492 -261 535 -255
rect 343 -306 352 -275
rect 492 -275 500 -261
rect 406 -306 414 -275
rect 343 -308 414 -306
rect 343 -309 415 -308
rect 190 -310 243 -309
rect 190 -322 216 -310
rect 242 -322 243 -310
rect 343 -314 440 -309
rect 190 -324 243 -322
rect 406 -318 440 -314
rect 232 -350 239 -334
rect 342 -342 391 -334
rect 249 -379 257 -359
rect 320 -376 328 -357
rect 342 -351 352 -342
rect 383 -349 391 -342
rect 406 -350 414 -318
rect 429 -323 440 -318
rect 515 -321 525 -288
rect 534 -321 1101 -320
rect 429 -333 470 -323
rect 515 -330 1101 -321
rect 515 -356 525 -330
rect 534 -331 1101 -330
rect 810 -332 868 -331
rect 225 -386 241 -379
rect 216 -387 219 -386
rect 249 -390 396 -379
rect 491 -383 500 -367
rect 1093 -373 1101 -331
rect 1400 -344 1423 -338
rect 1400 -354 1406 -344
rect 1564 -354 1570 -338
rect 1093 -374 1416 -373
rect 1093 -380 1409 -374
rect 1415 -380 1416 -374
rect 1419 -376 1425 -363
rect 1440 -376 1446 -363
rect 1419 -382 1446 -376
rect 1460 -376 1466 -363
rect 1479 -376 1485 -363
rect 1460 -382 1485 -376
rect 1498 -376 1504 -363
rect 1522 -376 1528 -363
rect 1498 -382 1528 -376
rect 491 -389 526 -383
rect 1541 -385 1547 -363
rect 1582 -384 1589 -362
rect 1582 -385 1596 -384
rect 1669 -385 1734 -384
rect 249 -391 404 -390
rect 1541 -391 1555 -385
rect 1582 -390 1734 -385
rect 249 -401 257 -391
rect 1541 -397 1547 -391
rect 232 -420 239 -410
rect 387 -414 395 -409
rect 582 -410 590 -402
rect 321 -415 445 -414
rect 450 -415 458 -410
rect 321 -420 458 -415
rect 321 -434 328 -420
rect 387 -421 458 -420
rect 387 -436 395 -421
rect 450 -437 458 -421
rect 547 -416 590 -410
rect 1419 -403 1547 -397
rect 1419 -415 1426 -403
rect 547 -430 555 -416
rect 1459 -415 1466 -403
rect 1498 -414 1505 -403
rect 343 -475 352 -444
rect 406 -475 414 -444
rect 343 -476 414 -475
rect 469 -476 477 -445
rect 343 -478 477 -476
rect 1400 -435 1406 -421
rect 1440 -435 1446 -421
rect 1540 -415 1547 -403
rect 1479 -435 1485 -422
rect 1582 -415 1589 -390
rect 1522 -435 1528 -422
rect 1400 -440 1528 -435
rect 1564 -438 1570 -421
rect 570 -476 580 -443
rect 585 -476 1158 -475
rect 1329 -476 1450 -475
rect 119 -480 197 -478
rect 136 -489 197 -480
rect 119 -491 197 -489
rect 343 -479 478 -478
rect 518 -479 525 -478
rect 343 -483 525 -479
rect 406 -487 525 -483
rect 469 -488 525 -487
rect 570 -484 1450 -476
rect 570 -485 1158 -484
rect 1329 -485 1450 -484
rect 234 -512 241 -497
rect 342 -511 391 -503
rect 82 -548 243 -541
rect 251 -548 259 -521
rect 320 -544 328 -526
rect 342 -520 352 -511
rect 383 -518 391 -511
rect 406 -512 454 -504
rect 406 -519 414 -512
rect 446 -519 454 -512
rect 469 -520 477 -488
rect 570 -511 580 -485
rect 546 -538 555 -522
rect 546 -544 581 -538
rect 251 -559 396 -548
rect 251 -560 404 -559
rect 251 -563 259 -560
rect 234 -582 241 -572
rect 367 -573 375 -568
rect 301 -574 425 -573
rect 430 -574 438 -569
rect 602 -571 610 -563
rect 301 -575 438 -574
rect 301 -576 493 -575
rect 498 -576 506 -571
rect 301 -579 506 -576
rect 301 -593 308 -579
rect 367 -580 506 -579
rect 367 -595 375 -580
rect 430 -582 506 -580
rect 430 -596 438 -582
rect 184 -634 216 -633
rect 323 -634 332 -603
rect 498 -598 506 -582
rect 567 -577 610 -571
rect 567 -591 575 -577
rect 386 -634 394 -603
rect 184 -650 197 -634
rect 323 -635 394 -634
rect 449 -635 457 -604
rect 323 -637 457 -635
rect 517 -637 525 -606
rect 323 -638 458 -637
rect 473 -638 525 -637
rect 323 -639 525 -638
rect 590 -637 600 -604
rect 590 -638 1158 -637
rect 1329 -638 1497 -637
rect 323 -640 526 -639
rect 538 -640 545 -639
rect 323 -642 545 -640
rect 386 -646 545 -642
rect 449 -647 545 -646
rect 481 -648 545 -647
rect 517 -649 545 -648
rect 590 -645 1488 -638
rect 1495 -645 1497 -638
rect 590 -646 617 -645
rect 1139 -646 1399 -645
rect 233 -667 240 -651
rect 322 -670 371 -662
rect 211 -696 214 -695
rect 211 -702 242 -696
rect 197 -703 242 -702
rect 250 -698 258 -676
rect 250 -707 282 -698
rect 300 -703 308 -685
rect 322 -679 332 -670
rect 363 -677 371 -670
rect 386 -671 434 -663
rect 449 -665 457 -664
rect 386 -678 394 -671
rect 426 -678 434 -671
rect 448 -672 502 -665
rect 449 -679 457 -672
rect 481 -673 502 -672
rect 494 -680 502 -673
rect 517 -681 525 -649
rect 590 -672 600 -646
rect 566 -699 575 -683
rect 566 -705 601 -699
rect 250 -708 376 -707
rect 250 -718 258 -708
rect 274 -718 376 -708
rect 975 -710 1115 -709
rect 975 -712 1099 -710
rect 275 -719 384 -718
rect 542 -721 1099 -712
rect 1114 -721 1115 -710
rect 542 -722 1115 -721
rect 233 -737 240 -727
rect 572 -763 1127 -761
rect 572 -773 574 -763
rect 583 -773 1127 -763
rect 572 -774 1142 -773
rect 376 -792 384 -787
rect 310 -793 434 -792
rect 439 -793 447 -788
rect 310 -794 447 -793
rect 310 -795 502 -794
rect 507 -795 515 -790
rect 672 -791 680 -783
rect 566 -795 574 -791
rect 310 -798 574 -795
rect 310 -812 317 -798
rect 376 -799 574 -798
rect 376 -814 384 -799
rect 439 -801 574 -799
rect 439 -815 447 -801
rect 505 -802 574 -801
rect 332 -853 341 -822
rect 507 -817 515 -802
rect 395 -853 403 -822
rect 332 -854 403 -853
rect 458 -854 466 -823
rect 566 -818 574 -802
rect 637 -797 680 -791
rect 637 -811 645 -797
rect 0 -856 210 -855
rect 332 -856 466 -854
rect 526 -856 534 -825
rect 0 -869 197 -856
rect 332 -857 467 -856
rect 482 -857 534 -856
rect 585 -857 593 -826
rect 332 -859 593 -857
rect 660 -857 670 -824
rect 674 -857 1158 -855
rect 1329 -857 1532 -855
rect 332 -860 594 -859
rect 606 -860 615 -859
rect 332 -861 615 -860
rect 395 -865 615 -861
rect 458 -866 615 -865
rect 490 -867 615 -866
rect 526 -868 615 -867
rect 585 -869 615 -868
rect 660 -865 1532 -857
rect 660 -866 687 -865
rect 0 -870 210 -869
rect 233 -899 240 -883
rect 331 -889 380 -881
rect 250 -925 258 -908
rect 283 -925 291 -924
rect 309 -925 317 -904
rect 331 -898 341 -889
rect 372 -896 380 -889
rect 395 -890 443 -882
rect 458 -884 466 -883
rect 395 -897 403 -890
rect 435 -897 443 -890
rect 457 -891 511 -884
rect 458 -898 466 -891
rect 490 -892 511 -891
rect 503 -899 511 -892
rect 526 -886 534 -885
rect 549 -886 570 -885
rect 526 -893 570 -886
rect 526 -900 534 -893
rect 562 -900 570 -893
rect 585 -901 593 -869
rect 660 -892 670 -866
rect 834 -867 881 -865
rect 1538 -865 1591 -855
rect 636 -919 645 -903
rect 636 -925 671 -919
rect -99 -928 216 -927
rect -99 -934 242 -928
rect -122 -935 242 -934
rect 250 -929 303 -925
rect 324 -926 335 -925
rect 324 -929 385 -926
rect 250 -936 385 -929
rect 250 -950 258 -936
rect 283 -937 385 -936
rect 846 -929 1113 -928
rect 846 -930 1097 -929
rect 631 -931 1097 -930
rect 551 -941 1097 -931
rect 233 -969 240 -959
<< m2contact >>
rect 40 1218 50 1231
rect 221 1421 234 1434
rect 204 1218 214 1231
rect 173 803 184 816
rect 155 488 161 495
rect 119 -489 136 -480
rect 174 -650 184 -633
rect -122 -934 -99 -927
<< metal2 >>
rect 18 1434 32 1435
rect 18 1422 221 1434
rect 18 1404 32 1422
rect -167 1390 32 1404
rect -124 541 -98 1390
rect 50 1218 204 1231
rect -122 -927 -99 541
rect 161 488 162 495
rect 155 357 162 488
rect -23 356 163 357
rect -34 348 163 356
rect -34 -480 -19 348
rect 155 0 162 348
rect -35 -489 119 -480
rect -34 -501 -19 -489
rect 174 -633 184 803
rect 174 -652 184 -650
rect -122 -936 -99 -934
<< labels >>
rlabel metal1 255 665 256 669 1 gnd
rlabel metal1 288 790 289 794 5 vdd
rlabel metal1 458 665 459 669 1 gnd
rlabel metal1 491 790 492 794 5 vdd
rlabel metal1 645 665 646 669 1 gnd
rlabel metal1 678 790 679 794 5 vdd
rlabel metal1 826 665 827 669 1 gnd
rlabel metal1 859 790 860 794 5 vdd
rlabel metal1 275 348 276 352 1 gnd
rlabel metal1 308 473 309 477 5 vdd
rlabel metal1 478 348 479 352 1 gnd
rlabel metal1 511 473 512 477 5 vdd
rlabel metal1 665 348 666 352 1 gnd
rlabel metal1 698 473 699 477 5 vdd
rlabel metal1 846 348 847 352 1 gnd
rlabel metal1 879 473 880 477 5 vdd
rlabel metal1 273 57 274 61 1 gnd
rlabel metal1 306 182 307 186 5 vdd
rlabel metal1 476 57 477 61 1 gnd
rlabel metal1 509 182 510 186 5 vdd
rlabel metal1 663 57 664 61 1 gnd
rlabel metal1 696 182 697 186 5 vdd
rlabel metal1 844 57 845 61 1 gnd
rlabel metal1 877 182 878 186 5 vdd
rlabel metal1 1231 505 1232 509 5 vdd
rlabel metal1 1198 380 1199 384 1 gnd
rlabel metal1 1368 506 1369 510 5 vdd
rlabel metal1 1462 485 1465 488 1 vdd
rlabel metal1 1462 408 1466 410 1 gnd
rlabel polysilicon 208 836 210 837 1 a1
rlabel polysilicon 244 519 246 520 1 a2
rlabel polysilicon 228 229 230 230 1 a3
rlabel polysilicon 207 809 209 810 1 b1
rlabel polycontact 223 490 225 491 1 b2
rlabel polycontact 221 200 223 201 1 b3
rlabel metal1 975 766 978 769 1 vdd
rlabel metal1 975 689 979 691 1 gnd
rlabel metal1 1000 372 1004 374 1 gnd
rlabel metal1 1000 449 1003 452 1 vdd
rlabel metal1 1009 81 1013 83 1 gnd
rlabel metal1 1009 158 1012 161 1 vdd
rlabel metal1 973 981 977 983 1 gnd
rlabel metal1 973 1058 976 1061 1 vdd
rlabel polysilicon 193 1097 195 1098 1 b0
rlabel polysilicon 200 1123 202 1124 1 a0
rlabel metal1 853 1079 854 1083 5 vdd
rlabel metal1 820 954 821 958 1 gnd
rlabel metal1 672 1079 673 1083 5 vdd
rlabel metal1 639 954 640 958 1 gnd
rlabel metal1 485 1079 486 1083 5 vdd
rlabel metal1 452 954 453 958 1 gnd
rlabel metal1 282 1079 283 1083 5 vdd
rlabel metal1 249 954 250 958 1 gnd
rlabel metal1 719 1343 721 1345 1 gnd
rlabel metal1 709 1472 711 1474 5 vdd
rlabel metal1 402 1469 403 1473 5 vdd
rlabel metal1 369 1344 370 1348 1 gnd
rlabel metal1 649 1563 651 1565 1 gnd
rlabel metal1 639 1692 641 1694 5 vdd
rlabel metal1 360 1563 361 1567 1 gnd
rlabel metal1 393 1688 394 1692 5 vdd
rlabel metal1 619 1853 621 1855 5 vdd
rlabel metal1 629 1724 631 1726 1 gnd
rlabel metal1 288 1608 291 1611 1 vdd
rlabel metal1 288 1531 292 1533 1 gnd
rlabel metal1 287 1848 291 1850 1 gnd
rlabel metal1 287 1925 290 1928 1 vdd
rlabel metal1 380 1722 381 1726 1 gnd
rlabel metal1 413 1847 414 1851 5 vdd
rlabel metal1 289 1763 292 1766 1 vdd
rlabel metal1 289 1686 293 1688 1 gnd
rlabel metal1 288 1299 292 1301 1 gnd
rlabel metal1 288 1376 291 1379 1 vdd
rlabel metal1 1506 1833 1507 1835 1 gnd
rlabel metal1 1506 1923 1507 1925 5 vdd
rlabel metal1 1483 1874 1484 1875 1 out
rlabel metal1 1343 1829 1344 1830 1 gnd
rlabel metal1 1344 1925 1345 1926 5 vdd
rlabel metal1 1512 442 1514 443 1 equal
rlabel metal1 564 2008 566 2010 5 vdd
rlabel metal1 574 1879 576 1881 1 gnd
rlabel metal1 413 2016 414 2020 5 vdd
rlabel metal1 380 1891 381 1895 1 gnd
rlabel metal1 1583 1878 1585 1879 1 agb
rlabel metal1 665 -923 667 -921 1 gnd
rlabel metal1 655 -794 657 -792 5 vdd
rlabel metal1 348 -797 349 -793 5 vdd
rlabel metal1 315 -922 316 -918 1 gnd
rlabel metal1 595 -703 597 -701 1 gnd
rlabel metal1 585 -574 587 -572 5 vdd
rlabel metal1 306 -703 307 -699 1 gnd
rlabel metal1 339 -578 340 -574 5 vdd
rlabel metal1 565 -413 567 -411 5 vdd
rlabel metal1 575 -542 577 -540 1 gnd
rlabel metal1 234 -658 237 -655 1 vdd
rlabel metal1 234 -735 238 -733 1 gnd
rlabel metal1 233 -418 237 -416 1 gnd
rlabel metal1 233 -341 236 -338 1 vdd
rlabel metal1 326 -544 327 -540 1 gnd
rlabel metal1 359 -419 360 -415 5 vdd
rlabel metal1 235 -503 238 -500 1 vdd
rlabel metal1 235 -580 239 -578 1 gnd
rlabel metal1 234 -967 238 -965 1 gnd
rlabel metal1 234 -890 237 -887 1 vdd
rlabel metal1 510 -258 512 -256 5 vdd
rlabel metal1 520 -387 522 -385 1 gnd
rlabel metal1 359 -250 360 -246 5 vdd
rlabel metal1 326 -375 327 -371 1 gnd
rlabel metal1 1404 -341 1405 -340 5 vdd
rlabel metal1 1403 -437 1404 -436 1 gnd
rlabel metal1 1566 -343 1567 -341 5 vdd
rlabel metal1 1566 -433 1567 -431 1 gnd
rlabel metal1 1643 -388 1644 -386 1 bga
<< end >>
